module master_control (
  clk,
  rst,
  mastertrig,
  hold_all_in,
  hold_buf_2,
  hold_buf_1,
  hold_buf_0,
  in_ctrl_buf_2,
  in_ctrl_buf_1,
  in_ctrl_buf_0,
  pos_hold_ctrl,
  Shuf_Ctrl_0,
  Shuf_Ctrl_1,
  Shuf_Ctrl_2,
  Shuf_Ctrl_3,
  Shuf_Ctrl_4,
  Shuf_Ctrl_5,
  Shuf_Ctrl_6,
  Shuf_Ctrl_7,
  Type_Sel_0,
  Type_Sel_1,
  Type_Sel_2,
  Type_Sel_3,
  Type_Sel_4,
  Type_Sel_5,
  Type_Sel_6,
  Type_Sel_7,
  Bypass_Sel_0,
  Bypass_Sel_1,
  Bypass_Sel_2,
  Bypass_Sel_3,
  Bypass_Sel_4,
  Bypass_Sel_5,
  Bypass_Sel_6,
  Bypass_Sel_7,
  DeShuf_Ctrl_0,
  DeShuf_Ctrl_1,
  DeShuf_Ctrl_2,
  DeShuf_Ctrl_3,
  DeShuf_Ctrl_4,
  DeShuf_Ctrl_5,
  DeShuf_Ctrl_6,
  DeShuf_Ctrl_7,
  Bypass_EN_0,
  Bypass_EN_1,
  Bypass_EN_2,
  Bypass_EN_3,
  Bypass_EN_4,
  Bypass_EN_5,
  Bypass_EN_6,
  Bypass_EN_7,
  Hold_Ctrl_0,
  Hold_Ctrl_1,
  Hold_Ctrl_2,
  Hold_Ctrl_3,
  Hold_Ctrl_4,
  Hold_Ctrl_5,
  Hold_Ctrl_6,
  Hold_Ctrl_7,
  DFF_Ctrl_0,
  DFF_Ctrl_1,
  DFF_Ctrl_2,
  DFF_Ctrl_3,
  DFF_Ctrl_4,
  DFF_Ctrl_5,
  DFF_Ctrl_6,
  DFF_Ctrl_7,
  hold_seg_0,
  hold_seg_1,
  hold_seg_2,
  hold_seg_3,
  hold_seg_4,
  hold_seg_5,
  hold_seg_6,
  hold_seg_7,
  in_ctrl_all_cb,
  hold_all_out,
  in_ctrl_all_out,
  counter_en
  );
  
  input                   clk;
  input                   rst;
  input                   mastertrig;
  output                  hold_all_in;
  output                  hold_buf_2;
  output                  hold_buf_1;
  output                  hold_buf_0;
  output                  in_ctrl_buf_2;
  output                  in_ctrl_buf_1;
  output                  in_ctrl_buf_0;
  output                  pos_hold_ctrl;
  output  [2:0]           Shuf_Ctrl_0;
  output  [2:0]           Shuf_Ctrl_1;
  output  [2:0]           Shuf_Ctrl_2;
  output  [2:0]           Shuf_Ctrl_3;
  output  [2:0]           Shuf_Ctrl_4;
  output  [2:0]           Shuf_Ctrl_5;
  output  [2:0]           Shuf_Ctrl_6;
  output  [2:0]           Shuf_Ctrl_7;
  output  [2:0]           Type_Sel_0;
  output  [2:0]           Type_Sel_1;
  output  [2:0]           Type_Sel_2;
  output  [2:0]           Type_Sel_3;
  output  [2:0]           Type_Sel_4;
  output  [2:0]           Type_Sel_5;
  output  [2:0]           Type_Sel_6;
  output  [2:0]           Type_Sel_7;
  output  [2:0]           Bypass_Sel_0;
  output  [2:0]           Bypass_Sel_1;
  output  [2:0]           Bypass_Sel_2;
  output  [2:0]           Bypass_Sel_3;
  output  [2:0]           Bypass_Sel_4;
  output  [2:0]           Bypass_Sel_5;
  output  [2:0]           Bypass_Sel_6;
  output  [2:0]           Bypass_Sel_7;
  output  [2:0]           DeShuf_Ctrl_0;
  output  [2:0]           DeShuf_Ctrl_1;
  output  [2:0]           DeShuf_Ctrl_2;
  output  [2:0]           DeShuf_Ctrl_3;
  output  [2:0]           DeShuf_Ctrl_4;
  output  [2:0]           DeShuf_Ctrl_5;
  output  [2:0]           DeShuf_Ctrl_6;
  output  [2:0]           DeShuf_Ctrl_7;
  output                  Bypass_EN_0;
  output                  Bypass_EN_1;
  output                  Bypass_EN_2;
  output                  Bypass_EN_3;
  output                  Bypass_EN_4;
  output                  Bypass_EN_5;
  output                  Bypass_EN_6;
  output                  Bypass_EN_7;
  output                  Hold_Ctrl_0;
  output                  Hold_Ctrl_1;
  output                  Hold_Ctrl_2;
  output                  Hold_Ctrl_3;
  output                  Hold_Ctrl_4;
  output                  Hold_Ctrl_5;
  output                  Hold_Ctrl_6;
  output                  Hold_Ctrl_7;
  output                  DFF_Ctrl_0;
  output                  DFF_Ctrl_1;
  output                  DFF_Ctrl_2;
  output                  DFF_Ctrl_3;
  output                  DFF_Ctrl_4;
  output                  DFF_Ctrl_5;
  output                  DFF_Ctrl_6;
  output                  DFF_Ctrl_7;
  output                  hold_seg_0;
  output                  hold_seg_1;
  output                  hold_seg_2;
  output                  hold_seg_3;
  output                  hold_seg_4;
  output                  hold_seg_5;
  output                  hold_seg_6;
  output                  hold_seg_7;
  output                  in_ctrl_all_cb;
  output                  hold_all_out;
  output                  in_ctrl_all_out;
  output                  counter_en;

  
  wire                    clk;
  wire                    rst;
  wire                    mastertrig;
  reg                     hold_all_in;
  reg                     hold_buf_2;
  reg                     hold_buf_1;
  reg                     hold_buf_0;
  reg                     in_ctrl_buf_2;
  reg                     in_ctrl_buf_1;
  reg                     in_ctrl_buf_0;
  reg                     pos_hold_ctrl;
  reg  [2:0]              Shuf_Ctrl_0;
  reg  [2:0]              Shuf_Ctrl_1;
  reg  [2:0]              Shuf_Ctrl_2;
  reg  [2:0]              Shuf_Ctrl_3;
  reg  [2:0]              Shuf_Ctrl_4;
  reg  [2:0]              Shuf_Ctrl_5;
  reg  [2:0]              Shuf_Ctrl_6;
  reg  [2:0]              Shuf_Ctrl_7;
  reg  [2:0]              Type_Sel_0;
  reg  [2:0]              Type_Sel_1;
  reg  [2:0]              Type_Sel_2;
  reg  [2:0]              Type_Sel_3;
  reg  [2:0]              Type_Sel_4;
  reg  [2:0]              Type_Sel_5;
  reg  [2:0]              Type_Sel_6;
  reg  [2:0]              Type_Sel_7;
  reg  [2:0]              Bypass_Sel_0;
  reg  [2:0]              Bypass_Sel_1;
  reg  [2:0]              Bypass_Sel_2;
  reg  [2:0]              Bypass_Sel_3;
  reg  [2:0]              Bypass_Sel_4;
  reg  [2:0]              Bypass_Sel_5;
  reg  [2:0]              Bypass_Sel_6;
  reg  [2:0]              Bypass_Sel_7;
  reg  [2:0]              DeShuf_Ctrl_0;
  reg  [2:0]              DeShuf_Ctrl_1;
  reg  [2:0]              DeShuf_Ctrl_2;
  reg  [2:0]              DeShuf_Ctrl_3;
  reg  [2:0]              DeShuf_Ctrl_4;
  reg  [2:0]              DeShuf_Ctrl_5;
  reg  [2:0]              DeShuf_Ctrl_6;
  reg  [2:0]              DeShuf_Ctrl_7;
  reg                     Bypass_EN_0;
  reg                     Bypass_EN_1;
  reg                     Bypass_EN_2;
  reg                     Bypass_EN_3;
  reg                     Bypass_EN_4;
  reg                     Bypass_EN_5;
  reg                     Bypass_EN_6;
  reg                     Bypass_EN_7;
  reg                     Hold_Ctrl_0;
  reg                     Hold_Ctrl_1;
  reg                     Hold_Ctrl_2;
  reg                     Hold_Ctrl_3;
  reg                     Hold_Ctrl_4;
  reg                     Hold_Ctrl_5;
  reg                     Hold_Ctrl_6;
  reg                     Hold_Ctrl_7;
  reg                     DFF_Ctrl_0;
  reg                     DFF_Ctrl_1;
  reg                     DFF_Ctrl_2;
  reg                     DFF_Ctrl_3;
  reg                     DFF_Ctrl_4;
  reg                     DFF_Ctrl_5;
  reg                     DFF_Ctrl_6;
  reg                     DFF_Ctrl_7;
  reg                     hold_seg_0;
  reg                     hold_seg_1;
  reg                     hold_seg_2;
  reg                     hold_seg_3;
  reg                     hold_seg_4;
  reg                     hold_seg_5;
  reg                     hold_seg_6;
  reg                     hold_seg_7;
  reg                     in_ctrl_all_cb;
  reg                     hold_all_out;
  reg                     in_ctrl_all_out;
  reg                     counter_en;
  
  localparam state_0  = 5'b00000;
  localparam state_1  = 5'b00001;
  localparam state_2  = 5'b00010;
  localparam state_3  = 5'b00011;
  localparam state_4  = 5'b00100;
  localparam state_5  = 5'b00101;
  localparam state_6  = 5'b00110;
  localparam state_7  = 5'b00111;
  localparam state_8  = 5'b01000;
  localparam state_9  = 5'b01001;
  localparam state_10 = 5'b01010;
  localparam state_11 = 5'b01011;
  localparam state_12 = 5'b01100;
  localparam state_13 = 5'b01101;
  localparam state_14 = 5'b01110;
  localparam state_15 = 5'b01111;
  localparam state_16 = 5'b10000;
  localparam state_17 = 5'b10001;
  localparam state_18 = 5'b10010;
  localparam state_19 = 5'b10011;
  localparam state_20 = 5'b10100;
  localparam state_21 = 5'b10101;
  localparam state_22 = 5'b10110;
  
  reg  [4:0] currentstate;
  
  always@(posedge clk)
    begin
      if(rst==1'b1)
        begin
          hold_all_in    <=  1'b0;
          hold_buf_2     <=  1'b1;
          hold_buf_1     <=  1'b1;
          hold_buf_0     <=  1'b1;
          in_ctrl_buf_2  <=  1'b0;
          in_ctrl_buf_1  <=  1'b0;
          in_ctrl_buf_0  <=  1'b0;
          pos_hold_ctrl  <=  1'b0;
          Shuf_Ctrl_0    <=  3'b000;
          Shuf_Ctrl_1    <=  3'b000;
          Shuf_Ctrl_2    <=  3'b000;
          Shuf_Ctrl_3    <=  3'b000;
          Shuf_Ctrl_4    <=  3'b000;
          Shuf_Ctrl_5    <=  3'b000;
          Shuf_Ctrl_6    <=  3'b000;
          Shuf_Ctrl_7    <=  3'b000;
          Type_Sel_0     <=  3'b000;
          Type_Sel_1     <=  3'b000;
          Type_Sel_2     <=  3'b000;
          Type_Sel_3     <=  3'b000;
          Type_Sel_4     <=  3'b000;
          Type_Sel_5     <=  3'b000;
          Type_Sel_6     <=  3'b000;
          Type_Sel_7     <=  3'b000;
          Bypass_Sel_0   <=  3'b000;
          Bypass_Sel_1   <=  3'b000;
          Bypass_Sel_2   <=  3'b000;
          Bypass_Sel_3   <=  3'b000;
          Bypass_Sel_4   <=  3'b000;
          Bypass_Sel_5   <=  3'b000;
          Bypass_Sel_6   <=  3'b000;
          Bypass_Sel_7   <=  3'b000;
          DeShuf_Ctrl_0  <=  3'b000;
          DeShuf_Ctrl_1  <=  3'b000;
          DeShuf_Ctrl_2  <=  3'b000;
          DeShuf_Ctrl_3  <=  3'b000;
          DeShuf_Ctrl_4  <=  3'b000;
          DeShuf_Ctrl_5  <=  3'b000;
          DeShuf_Ctrl_6  <=  3'b000;
          DeShuf_Ctrl_7  <=  3'b000;
          Bypass_EN_0    <=  1'b1;
          Bypass_EN_1    <=  1'b1;
          Bypass_EN_2    <=  1'b1;
          Bypass_EN_3    <=  1'b1;
          Bypass_EN_4    <=  1'b1;
          Bypass_EN_5    <=  1'b1;
          Bypass_EN_6    <=  1'b1;
          Bypass_EN_7    <=  1'b1;
          Hold_Ctrl_0    <=  1'b0;
          Hold_Ctrl_1    <=  1'b0;
          Hold_Ctrl_2    <=  1'b0;
          Hold_Ctrl_3    <=  1'b0;
          Hold_Ctrl_4    <=  1'b0;
          Hold_Ctrl_5    <=  1'b0;
          Hold_Ctrl_6    <=  1'b0;
          Hold_Ctrl_7    <=  1'b0;
          DFF_Ctrl_0     <=  1'b0;
          DFF_Ctrl_1     <=  1'b0;
          DFF_Ctrl_2     <=  1'b0;
          DFF_Ctrl_3     <=  1'b0;
          DFF_Ctrl_4     <=  1'b0;
          DFF_Ctrl_5     <=  1'b0;
          DFF_Ctrl_6     <=  1'b0;
          DFF_Ctrl_7     <=  1'b0;
          hold_seg_0     <=  1'b1;
          hold_seg_1     <=  1'b1;
          hold_seg_2     <=  1'b1;
          hold_seg_3     <=  1'b1;
          hold_seg_4     <=  1'b1;
          hold_seg_5     <=  1'b1;
          hold_seg_6     <=  1'b1;
          hold_seg_7     <=  1'b1;
          in_ctrl_all_cb <=  1'b1;
          hold_all_out   <=  1'b0;
          in_ctrl_all_out<=  1'b0;
          counter_en     <=  1'b0;	
          currentstate   <= state_0;          
        end
      else
        begin
          case(currentstate)
              state_0:
                begin
                  hold_all_in    <=  1'b0;
                  hold_buf_2     <=  1'b1;
                  hold_buf_1     <=  1'b1;
                  hold_buf_0     <=  1'b1;
                  in_ctrl_buf_2  <=  1'b0;
                  in_ctrl_buf_1  <=  1'b0;
                  in_ctrl_buf_0  <=  1'b0;
                  pos_hold_ctrl  <=  1'b0;
                  Shuf_Ctrl_0    <=  3'b000;
                  Shuf_Ctrl_1    <=  3'b000;
                  Shuf_Ctrl_2    <=  3'b000;
                  Shuf_Ctrl_3    <=  3'b000;
                  Shuf_Ctrl_4    <=  3'b000;
                  Shuf_Ctrl_5    <=  3'b000;
                  Shuf_Ctrl_6    <=  3'b000;
                  Shuf_Ctrl_7    <=  3'b000;
                  Type_Sel_0     <=  3'b000;
                  Type_Sel_1     <=  3'b000;
                  Type_Sel_2     <=  3'b000;
                  Type_Sel_3     <=  3'b000;
                  Type_Sel_4     <=  3'b000;
                  Type_Sel_5     <=  3'b000;
                  Type_Sel_6     <=  3'b000;
                  Type_Sel_7     <=  3'b000;
                  Bypass_Sel_0   <=  3'b000;
                  Bypass_Sel_1   <=  3'b000;
                  Bypass_Sel_2   <=  3'b000;
                  Bypass_Sel_3   <=  3'b000;
                  Bypass_Sel_4   <=  3'b000;
                  Bypass_Sel_5   <=  3'b000;
                  Bypass_Sel_6   <=  3'b000;
                  Bypass_Sel_7   <=  3'b000;
                  DeShuf_Ctrl_0  <=  3'b000;
                  DeShuf_Ctrl_1  <=  3'b000;
                  DeShuf_Ctrl_2  <=  3'b000;
                  DeShuf_Ctrl_3  <=  3'b000;
                  DeShuf_Ctrl_4  <=  3'b000;
                  DeShuf_Ctrl_5  <=  3'b000;
                  DeShuf_Ctrl_6  <=  3'b000;
                  DeShuf_Ctrl_7  <=  3'b000;
                  Bypass_EN_0    <=  1'b1;
                  Bypass_EN_1    <=  1'b1;
                  Bypass_EN_2    <=  1'b1;
                  Bypass_EN_3    <=  1'b1;
                  Bypass_EN_4    <=  1'b1;
                  Bypass_EN_5    <=  1'b1;
                  Bypass_EN_6    <=  1'b1;
                  Bypass_EN_7    <=  1'b1;
                  Hold_Ctrl_0    <=  1'b0;
                  Hold_Ctrl_1    <=  1'b0;
                  Hold_Ctrl_2    <=  1'b0;
                  Hold_Ctrl_3    <=  1'b0;
                  Hold_Ctrl_4    <=  1'b0;
                  Hold_Ctrl_5    <=  1'b0;
                  Hold_Ctrl_6    <=  1'b0;
                  Hold_Ctrl_7    <=  1'b0;
                  DFF_Ctrl_0     <=  1'b0;
                  DFF_Ctrl_1     <=  1'b0;
                  DFF_Ctrl_2     <=  1'b0;
                  DFF_Ctrl_3     <=  1'b0;
                  DFF_Ctrl_4     <=  1'b0;
                  DFF_Ctrl_5     <=  1'b0;
                  DFF_Ctrl_6     <=  1'b0;
                  DFF_Ctrl_7     <=  1'b0;
                  hold_seg_0     <=  1'b1;
                  hold_seg_1     <=  1'b1;
                  hold_seg_2     <=  1'b1;
                  hold_seg_3     <=  1'b1;
                  hold_seg_4     <=  1'b1;
                  hold_seg_5     <=  1'b1;
                  hold_seg_6     <=  1'b1;
                  hold_seg_7     <=  1'b1;
                  in_ctrl_all_cb <=  1'b1;
                  hold_all_out   <=  1'b0;
                  in_ctrl_all_out<=  1'b0;
                  counter_en     <=  1'b0;		
                  if (mastertrig==1'b1)
                    begin
                      currentstate <= state_1;
                    end
                  else
                    begin
                      currentstate <= state_0;
                    end
                end
              state_1:
                begin
                  hold_all_in    <=  1'b0;
                  hold_buf_2     <=  1'b1;
                  hold_buf_1     <=  1'b1;
                  hold_buf_0     <=  1'b1;
                  in_ctrl_buf_2  <=  1'b0;
                  in_ctrl_buf_1  <=  1'b0;
                  in_ctrl_buf_0  <=  1'b0;
                  pos_hold_ctrl  <=  1'b0;
                  Shuf_Ctrl_0    <=  3'b000;
                  Shuf_Ctrl_1    <=  3'b000;
                  Shuf_Ctrl_2    <=  3'b000;
                  Shuf_Ctrl_3    <=  3'b000;
                  Shuf_Ctrl_4    <=  3'b000;
                  Shuf_Ctrl_5    <=  3'b000;
                  Shuf_Ctrl_6    <=  3'b000;
                  Shuf_Ctrl_7    <=  3'b000;
                  Type_Sel_0     <=  3'b000;
                  Type_Sel_1     <=  3'b000;
                  Type_Sel_2     <=  3'b000;
                  Type_Sel_3     <=  3'b000;
                  Type_Sel_4     <=  3'b000;
                  Type_Sel_5     <=  3'b000;
                  Type_Sel_6     <=  3'b000;
                  Type_Sel_7     <=  3'b000;
                  Bypass_Sel_0   <=  3'b000;
                  Bypass_Sel_1   <=  3'b000;
                  Bypass_Sel_2   <=  3'b000;
                  Bypass_Sel_3   <=  3'b000;
                  Bypass_Sel_4   <=  3'b000;
                  Bypass_Sel_5   <=  3'b000;
                  Bypass_Sel_6   <=  3'b000;
                  Bypass_Sel_7   <=  3'b000;
                  DeShuf_Ctrl_0  <=  3'b000;
                  DeShuf_Ctrl_1  <=  3'b000;
                  DeShuf_Ctrl_2  <=  3'b000;
                  DeShuf_Ctrl_3  <=  3'b000;
                  DeShuf_Ctrl_4  <=  3'b000;
                  DeShuf_Ctrl_5  <=  3'b000;
                  DeShuf_Ctrl_6  <=  3'b000;
                  DeShuf_Ctrl_7  <=  3'b000;
                  Bypass_EN_0    <=  1'b1;
                  Bypass_EN_1    <=  1'b1;
                  Bypass_EN_2    <=  1'b1;
                  Bypass_EN_3    <=  1'b1;
                  Bypass_EN_4    <=  1'b1;
                  Bypass_EN_5    <=  1'b1;
                  Bypass_EN_6    <=  1'b1;
                  Bypass_EN_7    <=  1'b1;
                  Hold_Ctrl_0    <=  1'b0;
                  Hold_Ctrl_1    <=  1'b0;
                  Hold_Ctrl_2    <=  1'b0;
                  Hold_Ctrl_3    <=  1'b0;
                  Hold_Ctrl_4    <=  1'b0;
                  Hold_Ctrl_5    <=  1'b0;
                  Hold_Ctrl_6    <=  1'b0;
                  Hold_Ctrl_7    <=  1'b0;
                  DFF_Ctrl_0     <=  1'b0;
                  DFF_Ctrl_1     <=  1'b0;
                  DFF_Ctrl_2     <=  1'b0;
                  DFF_Ctrl_3     <=  1'b0;
                  DFF_Ctrl_4     <=  1'b0;
                  DFF_Ctrl_5     <=  1'b0;
                  DFF_Ctrl_6     <=  1'b0;
                  DFF_Ctrl_7     <=  1'b0;
                  hold_seg_0     <=  1'b0;
                  hold_seg_1     <=  1'b1;
                  hold_seg_2     <=  1'b1;
                  hold_seg_3     <=  1'b1;
                  hold_seg_4     <=  1'b1;
                  hold_seg_5     <=  1'b1;
                  hold_seg_6     <=  1'b1;
                  hold_seg_7     <=  1'b1;
                  in_ctrl_all_cb <=  1'b1;
                  hold_all_out   <=  1'b0;
                  in_ctrl_all_out<=  1'b0;
                  counter_en     <=  1'b0;
                  currentstate   <= state_2;
                end
              state_2:
                begin
                  hold_all_in    <=  1'b0;
                  hold_buf_2     <=  1'b1;
                  hold_buf_1     <=  1'b1;
                  hold_buf_0     <=  1'b1;
                  in_ctrl_buf_2  <=  1'b0;
                  in_ctrl_buf_1  <=  1'b0;
                  in_ctrl_buf_0  <=  1'b0;
                  pos_hold_ctrl  <=  1'b0;
                  Shuf_Ctrl_0    <=  3'b001;
                  Shuf_Ctrl_1    <=  3'b010;
                  Shuf_Ctrl_2    <=  3'b011;
                  Shuf_Ctrl_3    <=  3'b100;
                  Shuf_Ctrl_4    <=  3'b101;
                  Shuf_Ctrl_5    <=  3'b110;
                  Shuf_Ctrl_6    <=  3'b111;
                  Shuf_Ctrl_7    <=  3'b000;
                  Type_Sel_0     <=  3'b001;
                  Type_Sel_1     <=  3'b001;
                  Type_Sel_2     <=  3'b001;
                  Type_Sel_3     <=  3'b001;
                  Type_Sel_4     <=  3'b001;
                  Type_Sel_5     <=  3'b001;
                  Type_Sel_6     <=  3'b001;
                  Type_Sel_7     <=  3'b001;
                  Bypass_Sel_0   <=  3'b000;
                  Bypass_Sel_1   <=  3'b000;
                  Bypass_Sel_2   <=  3'b000;
                  Bypass_Sel_3   <=  3'b000;
                  Bypass_Sel_4   <=  3'b000;
                  Bypass_Sel_5   <=  3'b000;
                  Bypass_Sel_6   <=  3'b000;
                  Bypass_Sel_7   <=  3'b000;
                  DeShuf_Ctrl_0  <=  3'b000;
                  DeShuf_Ctrl_1  <=  3'b000;
                  DeShuf_Ctrl_2  <=  3'b001;
                  DeShuf_Ctrl_3  <=  3'b010;
                  DeShuf_Ctrl_4  <=  3'b011;
                  DeShuf_Ctrl_5  <=  3'b100;
                  DeShuf_Ctrl_6  <=  3'b101;
                  DeShuf_Ctrl_7  <=  3'b110;
                  Bypass_EN_0    <=  1'b1;
                  Bypass_EN_1    <=  1'b0;
                  Bypass_EN_2    <=  1'b0;
                  Bypass_EN_3    <=  1'b0;
                  Bypass_EN_4    <=  1'b0;
                  Bypass_EN_5    <=  1'b0;
                  Bypass_EN_6    <=  1'b0;
                  Bypass_EN_7    <=  1'b0;
                  Hold_Ctrl_0    <=  1'b0;
                  Hold_Ctrl_1    <=  1'b0;
                  Hold_Ctrl_2    <=  1'b0;
                  Hold_Ctrl_3    <=  1'b0;
                  Hold_Ctrl_4    <=  1'b0;
                  Hold_Ctrl_5    <=  1'b0;
                  Hold_Ctrl_6    <=  1'b0;
                  Hold_Ctrl_7    <=  1'b0;
                  DFF_Ctrl_0     <=  1'b0;
                  DFF_Ctrl_1     <=  1'b0;
                  DFF_Ctrl_2     <=  1'b0;
                  DFF_Ctrl_3     <=  1'b0;
                  DFF_Ctrl_4     <=  1'b0;
                  DFF_Ctrl_5     <=  1'b0;
                  DFF_Ctrl_6     <=  1'b0;
                  DFF_Ctrl_7     <=  1'b0;
                  hold_seg_0     <=  1'b1;
                  hold_seg_1     <=  1'b0;
                  hold_seg_2     <=  1'b1;
                  hold_seg_3     <=  1'b1;
                  hold_seg_4     <=  1'b1;
                  hold_seg_5     <=  1'b1;
                  hold_seg_6     <=  1'b1;
                  hold_seg_7     <=  1'b1;
                  in_ctrl_all_cb <=  1'b1;
                  hold_all_out   <=  1'b0;
                  in_ctrl_all_out<=  1'b0;
                  counter_en     <=  1'b0;
                  currentstate   <= state_3;
                end
              state_3:
                begin
                  hold_all_in    <=  1'b1;
                  hold_buf_2     <=  1'b1;
                  hold_buf_1     <=  1'b1;
                  hold_buf_0     <=  1'b0;
                  in_ctrl_buf_2  <=  1'b0;
                  in_ctrl_buf_1  <=  1'b0;
                  in_ctrl_buf_0  <=  1'b1;
                  pos_hold_ctrl  <=  1'b1;
                  Shuf_Ctrl_0    <=  3'b000;
                  Shuf_Ctrl_1    <=  3'b001;
                  Shuf_Ctrl_2    <=  3'b000;
                  Shuf_Ctrl_3    <=  3'b010;
                  Shuf_Ctrl_4    <=  3'b000;
                  Shuf_Ctrl_5    <=  3'b011;
                  Shuf_Ctrl_6    <=  3'b000;
                  Shuf_Ctrl_7    <=  3'b100;
                  Type_Sel_0     <=  3'b000;
                  Type_Sel_1     <=  3'b001;
                  Type_Sel_2     <=  3'b000;
                  Type_Sel_3     <=  3'b001;
                  Type_Sel_4     <=  3'b000;
                  Type_Sel_5     <=  3'b001;
                  Type_Sel_6     <=  3'b000;
                  Type_Sel_7     <=  3'b001;
                  Bypass_Sel_0   <=  3'b000;
                  Bypass_Sel_1   <=  3'b000;
                  Bypass_Sel_2   <=  3'b000;
                  Bypass_Sel_3   <=  3'b000;
                  Bypass_Sel_4   <=  3'b000;
                  Bypass_Sel_5   <=  3'b000;
                  Bypass_Sel_6   <=  3'b000;
                  Bypass_Sel_7   <=  3'b000;
                  DeShuf_Ctrl_0  <=  3'b000;
                  DeShuf_Ctrl_1  <=  3'b001;
                  DeShuf_Ctrl_2  <=  3'b011;
                  DeShuf_Ctrl_3  <=  3'b101;
                  DeShuf_Ctrl_4  <=  3'b111;
                  DeShuf_Ctrl_5  <=  3'b000;
                  DeShuf_Ctrl_6  <=  3'b000;
                  DeShuf_Ctrl_7  <=  3'b000;
                  Bypass_EN_0    <=  1'b1;
                  Bypass_EN_1    <=  1'b0;
                  Bypass_EN_2    <=  1'b0;
                  Bypass_EN_3    <=  1'b0;
                  Bypass_EN_4    <=  1'b0;
                  Bypass_EN_5    <=  1'b0;
                  Bypass_EN_6    <=  1'b0;
                  Bypass_EN_7    <=  1'b0;
                  Hold_Ctrl_0    <=  1'b0;
                  Hold_Ctrl_1    <=  1'b0;
                  Hold_Ctrl_2    <=  1'b0;
                  Hold_Ctrl_3    <=  1'b0;
                  Hold_Ctrl_4    <=  1'b0;
                  Hold_Ctrl_5    <=  1'b0;
                  Hold_Ctrl_6    <=  1'b0;
                  Hold_Ctrl_7    <=  1'b0;
                  DFF_Ctrl_0     <=  1'b0;
                  DFF_Ctrl_1     <=  1'b0;
                  DFF_Ctrl_2     <=  1'b0;
                  DFF_Ctrl_3     <=  1'b0;
                  DFF_Ctrl_4     <=  1'b0;
                  DFF_Ctrl_5     <=  1'b0;
                  DFF_Ctrl_6     <=  1'b0;
                  DFF_Ctrl_7     <=  1'b0;
                  hold_seg_0     <=  1'b1;
                  hold_seg_1     <=  1'b1;
                  hold_seg_2     <=  1'b1;
                  hold_seg_3     <=  1'b1;
                  hold_seg_4     <=  1'b1;
                  hold_seg_5     <=  1'b1;
                  hold_seg_6     <=  1'b1;
                  hold_seg_7     <=  1'b1;
                  in_ctrl_all_cb <=  1'b1;
                  hold_all_out   <=  1'b0;
                  in_ctrl_all_out<=  1'b0;
                  counter_en     <=  1'b0;
                  currentstate   <= state_4;
                end
              state_4:
                begin
                  hold_all_in    <=  1'b0;
                  hold_buf_2     <=  1'b1;
                  hold_buf_1     <=  1'b1;
                  hold_buf_0     <=  1'b0;
                  in_ctrl_buf_2  <=  1'b0;
                  in_ctrl_buf_1  <=  1'b0;
                  in_ctrl_buf_0  <=  1'b1;
                  pos_hold_ctrl  <=  1'b1;
                  Shuf_Ctrl_0    <=  3'b000;
                  Shuf_Ctrl_1    <=  3'b111;
                  Shuf_Ctrl_2    <=  3'b000;
                  Shuf_Ctrl_3    <=  3'b110;
                  Shuf_Ctrl_4    <=  3'b000;
                  Shuf_Ctrl_5    <=  3'b101;
                  Shuf_Ctrl_6    <=  3'b000;
                  Shuf_Ctrl_7    <=  3'b000;
                  Type_Sel_0     <=  3'b000;
                  Type_Sel_1     <=  3'b101;
                  Type_Sel_2     <=  3'b000;
                  Type_Sel_3     <=  3'b101;
                  Type_Sel_4     <=  3'b000;
                  Type_Sel_5     <=  3'b101;
                  Type_Sel_6     <=  3'b000;
                  Type_Sel_7     <=  3'b000;
                  Bypass_Sel_0   <=  3'b000;
                  Bypass_Sel_1   <=  3'b000;
                  Bypass_Sel_2   <=  3'b000;
                  Bypass_Sel_3   <=  3'b000;
                  Bypass_Sel_4   <=  3'b000;
                  Bypass_Sel_5   <=  3'b000;
                  Bypass_Sel_6   <=  3'b000;
                  Bypass_Sel_7   <=  3'b000;
                  DeShuf_Ctrl_0  <=  3'b000;
                  DeShuf_Ctrl_1  <=  3'b000;
                  DeShuf_Ctrl_2  <=  3'b000;
                  DeShuf_Ctrl_3  <=  3'b000;
                  DeShuf_Ctrl_4  <=  3'b000;
                  DeShuf_Ctrl_5  <=  3'b101;
                  DeShuf_Ctrl_6  <=  3'b011;
                  DeShuf_Ctrl_7  <=  3'b001;
                  Bypass_EN_0    <=  1'b1;
                  Bypass_EN_1    <=  1'b0;
                  Bypass_EN_2    <=  1'b0;
                  Bypass_EN_3    <=  1'b0;
                  Bypass_EN_4    <=  1'b0;
                  Bypass_EN_5    <=  1'b0;
                  Bypass_EN_6    <=  1'b0;
                  Bypass_EN_7    <=  1'b0;
                  Hold_Ctrl_0    <=  1'b1;
                  Hold_Ctrl_1    <=  1'b1;
                  Hold_Ctrl_2    <=  1'b1;
                  Hold_Ctrl_3    <=  1'b1;
                  Hold_Ctrl_4    <=  1'b1;
                  Hold_Ctrl_5    <=  1'b0;
                  Hold_Ctrl_6    <=  1'b0;
                  Hold_Ctrl_7    <=  1'b0;
                  DFF_Ctrl_0     <=  1'b1;
                  DFF_Ctrl_1     <=  1'b1;
                  DFF_Ctrl_2     <=  1'b1;
                  DFF_Ctrl_3     <=  1'b1;
                  DFF_Ctrl_4     <=  1'b1;
                  DFF_Ctrl_5     <=  1'b0;
                  DFF_Ctrl_6     <=  1'b0;
                  DFF_Ctrl_7     <=  1'b0;
                  hold_seg_0     <=  1'b1;
                  hold_seg_1     <=  1'b1;
                  hold_seg_2     <=  1'b0;
                  hold_seg_3     <=  1'b1;
                  hold_seg_4     <=  1'b1;
                  hold_seg_5     <=  1'b1;
                  hold_seg_6     <=  1'b1;
                  hold_seg_7     <=  1'b1;
                  in_ctrl_all_cb <=  1'b1;
                  hold_all_out   <=  1'b0;
                  in_ctrl_all_out<=  1'b0;
                  counter_en     <=  1'b0;
                  currentstate   <= state_5;
                end
              state_5:
                begin
                  hold_all_in    <=  1'b0;
                  hold_buf_2     <=  1'b1;
                  hold_buf_1     <=  1'b1;
                  hold_buf_0     <=  1'b0;
                  in_ctrl_buf_2  <=  1'b0;
                  in_ctrl_buf_1  <=  1'b0;
                  in_ctrl_buf_0  <=  1'b1;
                  pos_hold_ctrl  <=  1'b1;
                  Shuf_Ctrl_0    <=  3'b101;
                  Shuf_Ctrl_1    <=  3'b110;
                  Shuf_Ctrl_2    <=  3'b001;
                  Shuf_Ctrl_3    <=  3'b100;
                  Shuf_Ctrl_4    <=  3'b111;
                  Shuf_Ctrl_5    <=  3'b010;
                  Shuf_Ctrl_6    <=  3'b011;
                  Shuf_Ctrl_7    <=  3'b000;
                  Type_Sel_0     <=  3'b101;
                  Type_Sel_1     <=  3'b111;
                  Type_Sel_2     <=  3'b001;
                  Type_Sel_3     <=  3'b101;
                  Type_Sel_4     <=  3'b111;
                  Type_Sel_5     <=  3'b001;
                  Type_Sel_6     <=  3'b101;
                  Type_Sel_7     <=  3'b000;
                  Bypass_Sel_0   <=  3'b000;
                  Bypass_Sel_1   <=  3'b000;
                  Bypass_Sel_2   <=  3'b000;
                  Bypass_Sel_3   <=  3'b000;
                  Bypass_Sel_4   <=  3'b000;
                  Bypass_Sel_5   <=  3'b000;
                  Bypass_Sel_6   <=  3'b000;
                  Bypass_Sel_7   <=  3'b000;
                  DeShuf_Ctrl_0  <=  3'b000;
                  DeShuf_Ctrl_1  <=  3'b010;
                  DeShuf_Ctrl_2  <=  3'b101;
                  DeShuf_Ctrl_3  <=  3'b110;
                  DeShuf_Ctrl_4  <=  3'b011;
                  DeShuf_Ctrl_5  <=  3'b000;
                  DeShuf_Ctrl_6  <=  3'b001;
                  DeShuf_Ctrl_7  <=  3'b100;
                  Bypass_EN_0    <=  1'b1;
                  Bypass_EN_1    <=  1'b0;
                  Bypass_EN_2    <=  1'b0;
                  Bypass_EN_3    <=  1'b0;
                  Bypass_EN_4    <=  1'b0;
                  Bypass_EN_5    <=  1'b0;
                  Bypass_EN_6    <=  1'b0;
                  Bypass_EN_7    <=  1'b0;
                  Hold_Ctrl_0    <=  1'b0;
                  Hold_Ctrl_1    <=  1'b0;
                  Hold_Ctrl_2    <=  1'b0;
                  Hold_Ctrl_3    <=  1'b0;
                  Hold_Ctrl_4    <=  1'b0;
                  Hold_Ctrl_5    <=  1'b0;
                  Hold_Ctrl_6    <=  1'b0;
                  Hold_Ctrl_7    <=  1'b0;
                  DFF_Ctrl_0     <=  1'b0;
                  DFF_Ctrl_1     <=  1'b0;
                  DFF_Ctrl_2     <=  1'b0;
                  DFF_Ctrl_3     <=  1'b0;
                  DFF_Ctrl_4     <=  1'b0;
                  DFF_Ctrl_5     <=  1'b0;
                  DFF_Ctrl_6     <=  1'b0;
                  DFF_Ctrl_7     <=  1'b0;
                  hold_seg_0     <=  1'b1;
                  hold_seg_1     <=  1'b1;
                  hold_seg_2     <=  1'b1;
                  hold_seg_3     <=  1'b0;
                  hold_seg_4     <=  1'b1;
                  hold_seg_5     <=  1'b1;
                  hold_seg_6     <=  1'b1;
                  hold_seg_7     <=  1'b1;
                  in_ctrl_all_cb <=  1'b1;
                  hold_all_out   <=  1'b0;
                  in_ctrl_all_out<=  1'b0;
                  counter_en     <=  1'b0;
                  currentstate   <= state_6;
                end
              state_6:
                begin
                  hold_all_in    <=  1'b1;
                  hold_buf_2     <=  1'b1;
                  hold_buf_1     <=  1'b0;
                  hold_buf_0     <=  1'b1;
                  in_ctrl_buf_2  <=  1'b0;
                  in_ctrl_buf_1  <=  1'b1;
                  in_ctrl_buf_0  <=  1'b0;
                  pos_hold_ctrl  <=  1'b1;
                  Shuf_Ctrl_0    <=  3'b000;
                  Shuf_Ctrl_1    <=  3'b000;
                  Shuf_Ctrl_2    <=  3'b000;
                  Shuf_Ctrl_3    <=  3'b001;
                  Shuf_Ctrl_4    <=  3'b000;
                  Shuf_Ctrl_5    <=  3'b000;
                  Shuf_Ctrl_6    <=  3'b000;
                  Shuf_Ctrl_7    <=  3'b010;
                  Type_Sel_0     <=  3'b000;
                  Type_Sel_1     <=  3'b000;
                  Type_Sel_2     <=  3'b000;
                  Type_Sel_3     <=  3'b001;
                  Type_Sel_4     <=  3'b000;
                  Type_Sel_5     <=  3'b000;
                  Type_Sel_6     <=  3'b000;
                  Type_Sel_7     <=  3'b001;
                  Bypass_Sel_0   <=  3'b000;
                  Bypass_Sel_1   <=  3'b000;
                  Bypass_Sel_2   <=  3'b000;
                  Bypass_Sel_3   <=  3'b000;
                  Bypass_Sel_4   <=  3'b101;
                  Bypass_Sel_5   <=  3'b000;
                  Bypass_Sel_6   <=  3'b000;
                  Bypass_Sel_7   <=  3'b000;
                  DeShuf_Ctrl_0  <=  3'b000;
                  DeShuf_Ctrl_1  <=  3'b011;
                  DeShuf_Ctrl_2  <=  3'b111;
                  DeShuf_Ctrl_3  <=  3'b000;
                  DeShuf_Ctrl_4  <=  3'b000;
                  DeShuf_Ctrl_5  <=  3'b000;
                  DeShuf_Ctrl_6  <=  3'b000;
                  DeShuf_Ctrl_7  <=  3'b000;
                  Bypass_EN_0    <=  1'b1;
                  Bypass_EN_1    <=  1'b0;
                  Bypass_EN_2    <=  1'b0;
                  Bypass_EN_3    <=  1'b0;
                  Bypass_EN_4    <=  1'b1;
                  Bypass_EN_5    <=  1'b0;
                  Bypass_EN_6    <=  1'b0;
                  Bypass_EN_7    <=  1'b0;
                  Hold_Ctrl_0    <=  1'b0;
                  Hold_Ctrl_1    <=  1'b0;
                  Hold_Ctrl_2    <=  1'b0;
                  Hold_Ctrl_3    <=  1'b0;
                  Hold_Ctrl_4    <=  1'b0;
                  Hold_Ctrl_5    <=  1'b0;
                  Hold_Ctrl_6    <=  1'b0;
                  Hold_Ctrl_7    <=  1'b0;
                  DFF_Ctrl_0     <=  1'b0;
                  DFF_Ctrl_1     <=  1'b0;
                  DFF_Ctrl_2     <=  1'b0;
                  DFF_Ctrl_3     <=  1'b0;
                  DFF_Ctrl_4     <=  1'b0;
                  DFF_Ctrl_5     <=  1'b0;
                  DFF_Ctrl_6     <=  1'b0;
                  DFF_Ctrl_7     <=  1'b0;
                  hold_seg_0     <=  1'b1;
                  hold_seg_1     <=  1'b1;
                  hold_seg_2     <=  1'b1;
                  hold_seg_3     <=  1'b1;
                  hold_seg_4     <=  1'b1;
                  hold_seg_5     <=  1'b1;
                  hold_seg_6     <=  1'b1;
                  hold_seg_7     <=  1'b1;
                  in_ctrl_all_cb <=  1'b1;
                  hold_all_out   <=  1'b0;
                  in_ctrl_all_out<=  1'b0;
                  counter_en     <=  1'b0;
                  currentstate   <= state_7;
                end
              state_7:
                begin
                  hold_all_in    <=  1'b1;
                  hold_buf_2     <=  1'b0;
                  hold_buf_1     <=  1'b1;
                  hold_buf_0     <=  1'b1;
                  in_ctrl_buf_2  <=  1'b1;
                  in_ctrl_buf_1  <=  1'b0;
                  in_ctrl_buf_0  <=  1'b0;
                  pos_hold_ctrl  <=  1'b1;
                  Shuf_Ctrl_0    <=  3'b000;
                  Shuf_Ctrl_1    <=  3'b000;
                  Shuf_Ctrl_2    <=  3'b000;
                  Shuf_Ctrl_3    <=  3'b011;
                  Shuf_Ctrl_4    <=  3'b000;
                  Shuf_Ctrl_5    <=  3'b000;
                  Shuf_Ctrl_6    <=  3'b000;
                  Shuf_Ctrl_7    <=  3'b000;
                  Type_Sel_0     <=  3'b000;
                  Type_Sel_1     <=  3'b000;
                  Type_Sel_2     <=  3'b000;
                  Type_Sel_3     <=  3'b101;
                  Type_Sel_4     <=  3'b000;
                  Type_Sel_5     <=  3'b000;
                  Type_Sel_6     <=  3'b000;
                  Type_Sel_7     <=  3'b000;
                  Bypass_Sel_0   <=  3'b000;
                  Bypass_Sel_1   <=  3'b000;
                  Bypass_Sel_2   <=  3'b000;
                  Bypass_Sel_3   <=  3'b000;
                  Bypass_Sel_4   <=  3'b000;
                  Bypass_Sel_5   <=  3'b000;
                  Bypass_Sel_6   <=  3'b000;
                  Bypass_Sel_7   <=  3'b000;
                  DeShuf_Ctrl_0  <=  3'b000;
                  DeShuf_Ctrl_1  <=  3'b000;
                  DeShuf_Ctrl_2  <=  3'b000;
                  DeShuf_Ctrl_3  <=  3'b011;
                  DeShuf_Ctrl_4  <=  3'b000;
                  DeShuf_Ctrl_5  <=  3'b000;
                  DeShuf_Ctrl_6  <=  3'b000;
                  DeShuf_Ctrl_7  <=  3'b000;
                  Bypass_EN_0    <=  1'b1;
                  Bypass_EN_1    <=  1'b0;
                  Bypass_EN_2    <=  1'b0;
                  Bypass_EN_3    <=  1'b0;
                  Bypass_EN_4    <=  1'b0;
                  Bypass_EN_5    <=  1'b0;
                  Bypass_EN_6    <=  1'b0;
                  Bypass_EN_7    <=  1'b0;
                  Hold_Ctrl_0    <=  1'b1;
                  Hold_Ctrl_1    <=  1'b1;
                  Hold_Ctrl_2    <=  1'b1;
                  Hold_Ctrl_3    <=  1'b0;
                  Hold_Ctrl_4    <=  1'b1;
                  Hold_Ctrl_5    <=  1'b0;
                  Hold_Ctrl_6    <=  1'b0;
                  Hold_Ctrl_7    <=  1'b0;
                  DFF_Ctrl_0     <=  1'b1;
                  DFF_Ctrl_1     <=  1'b1;
                  DFF_Ctrl_2     <=  1'b1;
                  DFF_Ctrl_3     <=  1'b0;
                  DFF_Ctrl_4     <=  1'b1;
                  DFF_Ctrl_5     <=  1'b0;
                  DFF_Ctrl_6     <=  1'b0;
                  DFF_Ctrl_7     <=  1'b0;
                  hold_seg_0     <=  1'b1;
                  hold_seg_1     <=  1'b1;
                  hold_seg_2     <=  1'b1;
                  hold_seg_3     <=  1'b1;
                  hold_seg_4     <=  1'b1;
                  hold_seg_5     <=  1'b1;
                  hold_seg_6     <=  1'b1;
                  hold_seg_7     <=  1'b1;
                  in_ctrl_all_cb <=  1'b1;
                  hold_all_out   <=  1'b0;
                  in_ctrl_all_out<=  1'b0;
                  counter_en     <=  1'b0;
                  currentstate   <= state_8;
                end
              state_8:
                begin
                  hold_all_in    <=  1'b1;
                  hold_buf_2     <=  1'b1;
                  hold_buf_1     <=  1'b1;
                  hold_buf_0     <=  1'b1;
                  in_ctrl_buf_2  <=  1'b0;
                  in_ctrl_buf_1  <=  1'b0;
                  in_ctrl_buf_0  <=  1'b0;
                  pos_hold_ctrl  <=  1'b1;
                  Shuf_Ctrl_0    <=  3'b000;
                  Shuf_Ctrl_1    <=  3'b000;
                  Shuf_Ctrl_2    <=  3'b000;
                  Shuf_Ctrl_3    <=  3'b101;
                  Shuf_Ctrl_4    <=  3'b000;
                  Shuf_Ctrl_5    <=  3'b000;
                  Shuf_Ctrl_6    <=  3'b000;
                  Shuf_Ctrl_7    <=  3'b110;
                  Type_Sel_0     <=  3'b000;
                  Type_Sel_1     <=  3'b000;
                  Type_Sel_2     <=  3'b000;
                  Type_Sel_3     <=  3'b111;
                  Type_Sel_4     <=  3'b000;
                  Type_Sel_5     <=  3'b000;
                  Type_Sel_6     <=  3'b000;
                  Type_Sel_7     <=  3'b111;
                  Bypass_Sel_0   <=  3'b000;
                  Bypass_Sel_1   <=  3'b000;
                  Bypass_Sel_2   <=  3'b000;
                  Bypass_Sel_3   <=  3'b000;
                  Bypass_Sel_4   <=  3'b000;
                  Bypass_Sel_5   <=  3'b000;
                  Bypass_Sel_6   <=  3'b000;
                  Bypass_Sel_7   <=  3'b000;
                  DeShuf_Ctrl_0  <=  3'b000;
                  DeShuf_Ctrl_1  <=  3'b000;
                  DeShuf_Ctrl_2  <=  3'b000;
                  DeShuf_Ctrl_3  <=  3'b000;
                  DeShuf_Ctrl_4  <=  3'b000;
                  DeShuf_Ctrl_5  <=  3'b011;
                  DeShuf_Ctrl_6  <=  3'b111;
                  DeShuf_Ctrl_7  <=  3'b000;
                  Bypass_EN_0    <=  1'b1;
                  Bypass_EN_1    <=  1'b0;
                  Bypass_EN_2    <=  1'b0;
                  Bypass_EN_3    <=  1'b0;
                  Bypass_EN_4    <=  1'b0;
                  Bypass_EN_5    <=  1'b0;
                  Bypass_EN_6    <=  1'b0;
                  Bypass_EN_7    <=  1'b0;
                  Hold_Ctrl_0    <=  1'b1;
                  Hold_Ctrl_1    <=  1'b1;
                  Hold_Ctrl_2    <=  1'b1;
                  Hold_Ctrl_3    <=  1'b1;
                  Hold_Ctrl_4    <=  1'b1;
                  Hold_Ctrl_5    <=  1'b0;
                  Hold_Ctrl_6    <=  1'b0;
                  Hold_Ctrl_7    <=  1'b0;
                  DFF_Ctrl_0     <=  1'b1;
                  DFF_Ctrl_1     <=  1'b1;
                  DFF_Ctrl_2     <=  1'b1;
                  DFF_Ctrl_3     <=  1'b1;
                  DFF_Ctrl_4     <=  1'b1;
                  DFF_Ctrl_5     <=  1'b0;
                  DFF_Ctrl_6     <=  1'b0;
                  DFF_Ctrl_7     <=  1'b0;
                  hold_seg_0     <=  1'b1;
                  hold_seg_1     <=  1'b1;
                  hold_seg_2     <=  1'b1;
                  hold_seg_3     <=  1'b1;
                  hold_seg_4     <=  1'b1;
                  hold_seg_5     <=  1'b1;
                  hold_seg_6     <=  1'b1;
                  hold_seg_7     <=  1'b1;
                  in_ctrl_all_cb <=  1'b1;
                  hold_all_out   <=  1'b0;
                  in_ctrl_all_out<=  1'b0;
                  counter_en     <=  1'b0;
                  currentstate   <= state_9;
                end
              state_9:
                begin
                  hold_all_in    <=  1'b0;
                  hold_buf_2     <=  1'b0;
                  hold_buf_1     <=  1'b0;
                  hold_buf_0     <=  1'b0;
                  in_ctrl_buf_2  <=  1'b0;
                  in_ctrl_buf_1  <=  1'b0;
                  in_ctrl_buf_0  <=  1'b0;
                  pos_hold_ctrl  <=  1'b1;
                  Shuf_Ctrl_0    <=  3'b000;
                  Shuf_Ctrl_1    <=  3'b000;
                  Shuf_Ctrl_2    <=  3'b000;
                  Shuf_Ctrl_3    <=  3'b111;
                  Shuf_Ctrl_4    <=  3'b000;
                  Shuf_Ctrl_5    <=  3'b000;
                  Shuf_Ctrl_6    <=  3'b000;
                  Shuf_Ctrl_7    <=  3'b000;
                  Type_Sel_0     <=  3'b000;
                  Type_Sel_1     <=  3'b000;
                  Type_Sel_2     <=  3'b000;
                  Type_Sel_3     <=  3'b011;
                  Type_Sel_4     <=  3'b000;
                  Type_Sel_5     <=  3'b000;
                  Type_Sel_6     <=  3'b000;
                  Type_Sel_7     <=  3'b000;
                  Bypass_Sel_0   <=  3'b000;
                  Bypass_Sel_1   <=  3'b000;
                  Bypass_Sel_2   <=  3'b000;
                  Bypass_Sel_3   <=  3'b000;
                  Bypass_Sel_4   <=  3'b000;
                  Bypass_Sel_5   <=  3'b000;
                  Bypass_Sel_6   <=  3'b000;
                  Bypass_Sel_7   <=  3'b000;
                  DeShuf_Ctrl_0  <=  3'b000;
                  DeShuf_Ctrl_1  <=  3'b000;
                  DeShuf_Ctrl_2  <=  3'b000;
                  DeShuf_Ctrl_3  <=  3'b000;
                  DeShuf_Ctrl_4  <=  3'b000;
                  DeShuf_Ctrl_5  <=  3'b000;
                  DeShuf_Ctrl_6  <=  3'b000;
                  DeShuf_Ctrl_7  <=  3'b011;
                  Bypass_EN_0    <=  1'b1;
                  Bypass_EN_1    <=  1'b0;
                  Bypass_EN_2    <=  1'b0;
                  Bypass_EN_3    <=  1'b0;
                  Bypass_EN_4    <=  1'b0;
                  Bypass_EN_5    <=  1'b0;
                  Bypass_EN_6    <=  1'b0;
                  Bypass_EN_7    <=  1'b0;
                  Hold_Ctrl_0    <=  1'b1;
                  Hold_Ctrl_1    <=  1'b1;
                  Hold_Ctrl_2    <=  1'b1;
                  Hold_Ctrl_3    <=  1'b1;
                  Hold_Ctrl_4    <=  1'b1;
                  Hold_Ctrl_5    <=  1'b1;
                  Hold_Ctrl_6    <=  1'b1;
                  Hold_Ctrl_7    <=  1'b0;
                  DFF_Ctrl_0     <=  1'b1;
                  DFF_Ctrl_1     <=  1'b1;
                  DFF_Ctrl_2     <=  1'b1;
                  DFF_Ctrl_3     <=  1'b1;
                  DFF_Ctrl_4     <=  1'b1;
                  DFF_Ctrl_5     <=  1'b1;
                  DFF_Ctrl_6     <=  1'b1;
                  DFF_Ctrl_7     <=  1'b0;
                  hold_seg_0     <=  1'b1;
                  hold_seg_1     <=  1'b1;
                  hold_seg_2     <=  1'b1;
                  hold_seg_3     <=  1'b1;
                  hold_seg_4     <=  1'b0;
                  hold_seg_5     <=  1'b1;
                  hold_seg_6     <=  1'b1;
                  hold_seg_7     <=  1'b1;
                  in_ctrl_all_cb <=  1'b1;
                  hold_all_out   <=  1'b0;
                  in_ctrl_all_out<=  1'b0;
                  counter_en     <=  1'b0;
                  currentstate   <= state_10;
                end
              state_10:
                begin
                  hold_all_in    <=  1'b0;
                  hold_buf_2     <=  1'b0;
                  hold_buf_1     <=  1'b0;
                  hold_buf_0     <=  1'b0;
                  in_ctrl_buf_2  <=  1'b0;
                  in_ctrl_buf_1  <=  1'b0;
                  in_ctrl_buf_0  <=  1'b0;
                  pos_hold_ctrl  <=  1'b1;
                  Shuf_Ctrl_0    <=  3'b011;
                  Shuf_Ctrl_1    <=  3'b110;
                  Shuf_Ctrl_2    <=  3'b111;
                  Shuf_Ctrl_3    <=  3'b100;
                  Shuf_Ctrl_4    <=  3'b001;
                  Shuf_Ctrl_5    <=  3'b010;
                  Shuf_Ctrl_6    <=  3'b101;
                  Shuf_Ctrl_7    <=  3'b000;
                  Type_Sel_0     <=  3'b101;
                  Type_Sel_1     <=  3'b011;
                  Type_Sel_2     <=  3'b010;
                  Type_Sel_3     <=  3'b111;
                  Type_Sel_4     <=  3'b001;
                  Type_Sel_5     <=  3'b101;
                  Type_Sel_6     <=  3'b011;
                  Type_Sel_7     <=  3'b000;
                  Bypass_Sel_0   <=  3'b000;
                  Bypass_Sel_1   <=  3'b000;
                  Bypass_Sel_2   <=  3'b000;
                  Bypass_Sel_3   <=  3'b000;
                  Bypass_Sel_4   <=  3'b000;
                  Bypass_Sel_5   <=  3'b000;
                  Bypass_Sel_6   <=  3'b000;
                  Bypass_Sel_7   <=  3'b000;
                  DeShuf_Ctrl_0  <=  3'b000;
                  DeShuf_Ctrl_1  <=  3'b100;
                  DeShuf_Ctrl_2  <=  3'b101;
                  DeShuf_Ctrl_3  <=  3'b000;
                  DeShuf_Ctrl_4  <=  3'b011;
                  DeShuf_Ctrl_5  <=  3'b110;
                  DeShuf_Ctrl_6  <=  3'b001;
                  DeShuf_Ctrl_7  <=  3'b010;
                  Bypass_EN_0    <=  1'b1;
                  Bypass_EN_1    <=  1'b0;
                  Bypass_EN_2    <=  1'b0;
                  Bypass_EN_3    <=  1'b0;
                  Bypass_EN_4    <=  1'b0;
                  Bypass_EN_5    <=  1'b0;
                  Bypass_EN_6    <=  1'b0;
                  Bypass_EN_7    <=  1'b0;
                  Hold_Ctrl_0    <=  1'b0;
                  Hold_Ctrl_1    <=  1'b0;
                  Hold_Ctrl_2    <=  1'b0;
                  Hold_Ctrl_3    <=  1'b0;
                  Hold_Ctrl_4    <=  1'b0;
                  Hold_Ctrl_5    <=  1'b0;
                  Hold_Ctrl_6    <=  1'b0;
                  Hold_Ctrl_7    <=  1'b0;
                  DFF_Ctrl_0     <=  1'b0;
                  DFF_Ctrl_1     <=  1'b0;
                  DFF_Ctrl_2     <=  1'b0;
                  DFF_Ctrl_3     <=  1'b0;
                  DFF_Ctrl_4     <=  1'b0;
                  DFF_Ctrl_5     <=  1'b0;
                  DFF_Ctrl_6     <=  1'b0;
                  DFF_Ctrl_7     <=  1'b0;
                  hold_seg_0     <=  1'b1;
                  hold_seg_1     <=  1'b1;
                  hold_seg_2     <=  1'b1;
                  hold_seg_3     <=  1'b1;
                  hold_seg_4     <=  1'b1;
                  hold_seg_5     <=  1'b0;
                  hold_seg_6     <=  1'b1;
                  hold_seg_7     <=  1'b1;
                  in_ctrl_all_cb <=  1'b1;
                  hold_all_out   <=  1'b0;
                  in_ctrl_all_out<=  1'b0;
                  counter_en     <=  1'b0;
                  currentstate   <= state_11;
                end
              state_11:
                begin
                  hold_all_in    <=  1'b1;
                  hold_buf_2     <=  1'b1;
                  hold_buf_1     <=  1'b1;
                  hold_buf_0     <=  1'b1;
                  in_ctrl_buf_2  <=  1'b0;
                  in_ctrl_buf_1  <=  1'b0;
                  in_ctrl_buf_0  <=  1'b0;
                  pos_hold_ctrl  <=  1'b1;
                  Shuf_Ctrl_0    <=  3'b000;
                  Shuf_Ctrl_1    <=  3'b011;
                  Shuf_Ctrl_2    <=  3'b000;
                  Shuf_Ctrl_3    <=  3'b010;
                  Shuf_Ctrl_4    <=  3'b000;
                  Shuf_Ctrl_5    <=  3'b001;
                  Shuf_Ctrl_6    <=  3'b000;
                  Shuf_Ctrl_7    <=  3'b100;
                  Type_Sel_0     <=  3'b000;
                  Type_Sel_1     <=  3'b111;
                  Type_Sel_2     <=  3'b000;
                  Type_Sel_3     <=  3'b101;
                  Type_Sel_4     <=  3'b000;
                  Type_Sel_5     <=  3'b001;
                  Type_Sel_6     <=  3'b000;
                  Type_Sel_7     <=  3'b111;
                  Bypass_Sel_0   <=  3'b000;
                  Bypass_Sel_1   <=  3'b000;
                  Bypass_Sel_2   <=  3'b000;
                  Bypass_Sel_3   <=  3'b000;
                  Bypass_Sel_4   <=  3'b000;
                  Bypass_Sel_5   <=  3'b000;
                  Bypass_Sel_6   <=  3'b000;
                  Bypass_Sel_7   <=  3'b000;
                  DeShuf_Ctrl_0  <=  3'b000;
                  DeShuf_Ctrl_1  <=  3'b101;
                  DeShuf_Ctrl_2  <=  3'b011;
                  DeShuf_Ctrl_3  <=  3'b001;
                  DeShuf_Ctrl_4  <=  3'b111;
                  DeShuf_Ctrl_5  <=  3'b000;
                  DeShuf_Ctrl_6  <=  3'b000;
                  DeShuf_Ctrl_7  <=  3'b000;
                  Bypass_EN_0    <=  1'b1;
                  Bypass_EN_1    <=  1'b0;
                  Bypass_EN_2    <=  1'b0;
                  Bypass_EN_3    <=  1'b0;
                  Bypass_EN_4    <=  1'b0;
                  Bypass_EN_5    <=  1'b0;
                  Bypass_EN_6    <=  1'b0;
                  Bypass_EN_7    <=  1'b0;
                  Hold_Ctrl_0    <=  1'b0;
                  Hold_Ctrl_1    <=  1'b0;
                  Hold_Ctrl_2    <=  1'b0;
                  Hold_Ctrl_3    <=  1'b0;
                  Hold_Ctrl_4    <=  1'b0;
                  Hold_Ctrl_5    <=  1'b0;
                  Hold_Ctrl_6    <=  1'b0;
                  Hold_Ctrl_7    <=  1'b0;
                  DFF_Ctrl_0     <=  1'b0;
                  DFF_Ctrl_1     <=  1'b0;
                  DFF_Ctrl_2     <=  1'b0;
                  DFF_Ctrl_3     <=  1'b0;
                  DFF_Ctrl_4     <=  1'b0;
                  DFF_Ctrl_5     <=  1'b0;
                  DFF_Ctrl_6     <=  1'b0;
                  DFF_Ctrl_7     <=  1'b0;
                  hold_seg_0     <=  1'b1;
                  hold_seg_1     <=  1'b1;
                  hold_seg_2     <=  1'b1;
                  hold_seg_3     <=  1'b1;
                  hold_seg_4     <=  1'b1;
                  hold_seg_5     <=  1'b1;
                  hold_seg_6     <=  1'b1;
                  hold_seg_7     <=  1'b1;
                  in_ctrl_all_cb <=  1'b1;
                  hold_all_out   <=  1'b0;
                  in_ctrl_all_out<=  1'b0;
                  counter_en     <=  1'b0;
                  currentstate   <= state_12;
                end
              state_12:
                begin
                  hold_all_in    <=  1'b0;
                  hold_buf_2     <=  1'b0;
                  hold_buf_1     <=  1'b0;
                  hold_buf_0     <=  1'b0;
                  in_ctrl_buf_2  <=  1'b0;
                  in_ctrl_buf_1  <=  1'b0;
                  in_ctrl_buf_0  <=  1'b0;
                  pos_hold_ctrl  <=  1'b1;
                  Shuf_Ctrl_0    <=  3'b000;
                  Shuf_Ctrl_1    <=  3'b101;
                  Shuf_Ctrl_2    <=  3'b000;
                  Shuf_Ctrl_3    <=  3'b110;
                  Shuf_Ctrl_4    <=  3'b000;
                  Shuf_Ctrl_5    <=  3'b111;
                  Shuf_Ctrl_6    <=  3'b000;
                  Shuf_Ctrl_7    <=  3'b000;
                  Type_Sel_0     <=  3'b000;
                  Type_Sel_1     <=  3'b011;
                  Type_Sel_2     <=  3'b000;
                  Type_Sel_3     <=  3'b010;
                  Type_Sel_4     <=  3'b000;
                  Type_Sel_5     <=  3'b110;
                  Type_Sel_6     <=  3'b000;
                  Type_Sel_7     <=  3'b000;
                  Bypass_Sel_0   <=  3'b000;
                  Bypass_Sel_1   <=  3'b000;
                  Bypass_Sel_2   <=  3'b000;
                  Bypass_Sel_3   <=  3'b000;
                  Bypass_Sel_4   <=  3'b000;
                  Bypass_Sel_5   <=  3'b000;
                  Bypass_Sel_6   <=  3'b000;
                  Bypass_Sel_7   <=  3'b000;
                  DeShuf_Ctrl_0  <=  3'b000;
                  DeShuf_Ctrl_1  <=  3'b000;
                  DeShuf_Ctrl_2  <=  3'b000;
                  DeShuf_Ctrl_3  <=  3'b000;
                  DeShuf_Ctrl_4  <=  3'b000;
                  DeShuf_Ctrl_5  <=  3'b001;
                  DeShuf_Ctrl_6  <=  3'b011;
                  DeShuf_Ctrl_7  <=  3'b101;
                  Bypass_EN_0    <=  1'b1;
                  Bypass_EN_1    <=  1'b0;
                  Bypass_EN_2    <=  1'b0;
                  Bypass_EN_3    <=  1'b0;
                  Bypass_EN_4    <=  1'b0;
                  Bypass_EN_5    <=  1'b0;
                  Bypass_EN_6    <=  1'b0;
                  Bypass_EN_7    <=  1'b0;
                  Hold_Ctrl_0    <=  1'b1;
                  Hold_Ctrl_1    <=  1'b1;
                  Hold_Ctrl_2    <=  1'b1;
                  Hold_Ctrl_3    <=  1'b1;
                  Hold_Ctrl_4    <=  1'b1;
                  Hold_Ctrl_5    <=  1'b0;
                  Hold_Ctrl_6    <=  1'b0;
                  Hold_Ctrl_7    <=  1'b0;
                  DFF_Ctrl_0     <=  1'b1;
                  DFF_Ctrl_1     <=  1'b1;
                  DFF_Ctrl_2     <=  1'b1;
                  DFF_Ctrl_3     <=  1'b1;
                  DFF_Ctrl_4     <=  1'b1;
                  DFF_Ctrl_5     <=  1'b0;
                  DFF_Ctrl_6     <=  1'b0;
                  DFF_Ctrl_7     <=  1'b0;
                  hold_seg_0     <=  1'b1;
                  hold_seg_1     <=  1'b1;
                  hold_seg_2     <=  1'b1;
                  hold_seg_3     <=  1'b1;
                  hold_seg_4     <=  1'b1;
                  hold_seg_5     <=  1'b1;
                  hold_seg_6     <=  1'b0;
                  hold_seg_7     <=  1'b1;
                  in_ctrl_all_cb <=  1'b1;
                  hold_all_out   <=  1'b0;
                  in_ctrl_all_out<=  1'b0;
                  counter_en     <=  1'b0;
                  currentstate   <= state_13;
                end
              state_13:
                begin
                  hold_all_in    <=  1'b0;
                  hold_buf_2     <=  1'b1;
                  hold_buf_1     <=  1'b1;
                  hold_buf_0     <=  1'b1;
                  in_ctrl_buf_2  <=  1'b0;
                  in_ctrl_buf_1  <=  1'b0;
                  in_ctrl_buf_0  <=  1'b0;
                  pos_hold_ctrl  <=  1'b0;
                  Shuf_Ctrl_0    <=  3'b111;
                  Shuf_Ctrl_1    <=  3'b010;
                  Shuf_Ctrl_2    <=  3'b101;
                  Shuf_Ctrl_3    <=  3'b100;
                  Shuf_Ctrl_4    <=  3'b011;
                  Shuf_Ctrl_5    <=  3'b110;
                  Shuf_Ctrl_6    <=  3'b001;
                  Shuf_Ctrl_7    <=  3'b000;
                  Type_Sel_0     <=  3'b100;
                  Type_Sel_1     <=  3'b101;
                  Type_Sel_2     <=  3'b010;
                  Type_Sel_3     <=  3'b011;
                  Type_Sel_4     <=  3'b111;
                  Type_Sel_5     <=  3'b110;
                  Type_Sel_6     <=  3'b001;
                  Type_Sel_7     <=  3'b000;
                  Bypass_Sel_0   <=  3'b000;
                  Bypass_Sel_1   <=  3'b000;
                  Bypass_Sel_2   <=  3'b000;
                  Bypass_Sel_3   <=  3'b000;
                  Bypass_Sel_4   <=  3'b000;
                  Bypass_Sel_5   <=  3'b000;
                  Bypass_Sel_6   <=  3'b000;
                  Bypass_Sel_7   <=  3'b000;
                  DeShuf_Ctrl_0  <=  3'b000;
                  DeShuf_Ctrl_1  <=  3'b110;
                  DeShuf_Ctrl_2  <=  3'b001;
                  DeShuf_Ctrl_3  <=  3'b100;
                  DeShuf_Ctrl_4  <=  3'b011;
                  DeShuf_Ctrl_5  <=  3'b010;
                  DeShuf_Ctrl_6  <=  3'b101;
                  DeShuf_Ctrl_7  <=  3'b000;
                  Bypass_EN_0    <=  1'b1;
                  Bypass_EN_1    <=  1'b0;
                  Bypass_EN_2    <=  1'b0;
                  Bypass_EN_3    <=  1'b0;
                  Bypass_EN_4    <=  1'b0;
                  Bypass_EN_5    <=  1'b0;
                  Bypass_EN_6    <=  1'b0;
                  Bypass_EN_7    <=  1'b0;
                  Hold_Ctrl_0    <=  1'b0;
                  Hold_Ctrl_1    <=  1'b0;
                  Hold_Ctrl_2    <=  1'b0;
                  Hold_Ctrl_3    <=  1'b0;
                  Hold_Ctrl_4    <=  1'b0;
                  Hold_Ctrl_5    <=  1'b0;
                  Hold_Ctrl_6    <=  1'b0;
                  Hold_Ctrl_7    <=  1'b0;
                  DFF_Ctrl_0     <=  1'b0;
                  DFF_Ctrl_1     <=  1'b0;
                  DFF_Ctrl_2     <=  1'b0;
                  DFF_Ctrl_3     <=  1'b0;
                  DFF_Ctrl_4     <=  1'b0;
                  DFF_Ctrl_5     <=  1'b0;
                  DFF_Ctrl_6     <=  1'b0;
                  DFF_Ctrl_7     <=  1'b0;
                  hold_seg_0     <=  1'b1;
                  hold_seg_1     <=  1'b1;
                  hold_seg_2     <=  1'b1;
                  hold_seg_3     <=  1'b1;
                  hold_seg_4     <=  1'b1;
                  hold_seg_5     <=  1'b1;
                  hold_seg_6     <=  1'b1;
                  hold_seg_7     <=  1'b0;
                  in_ctrl_all_cb <=  1'b1;
                  hold_all_out   <=  1'b0;
                  in_ctrl_all_out<=  1'b1;
                  counter_en     <=  1'b0;
                  currentstate   <= state_14;
                end
              state_14:
                begin
                  hold_all_in    <=  1'b0;
                  hold_buf_2     <=  1'b1;
                  hold_buf_1     <=  1'b1;
                  hold_buf_0     <=  1'b1;
                  in_ctrl_buf_2  <=  1'b0;
                  in_ctrl_buf_1  <=  1'b0;
                  in_ctrl_buf_0  <=  1'b0;
                  pos_hold_ctrl  <=  1'b0;
                  Shuf_Ctrl_0    <=  3'b000;
                  Shuf_Ctrl_1    <=  3'b000;
                  Shuf_Ctrl_2    <=  3'b000;
                  Shuf_Ctrl_3    <=  3'b000;
                  Shuf_Ctrl_4    <=  3'b000;
                  Shuf_Ctrl_5    <=  3'b000;
                  Shuf_Ctrl_6    <=  3'b000;
                  Shuf_Ctrl_7    <=  3'b000;
                  Type_Sel_0     <=  3'b000;
                  Type_Sel_1     <=  3'b000;
                  Type_Sel_2     <=  3'b000;
                  Type_Sel_3     <=  3'b000;
                  Type_Sel_4     <=  3'b000;
                  Type_Sel_5     <=  3'b000;
                  Type_Sel_6     <=  3'b000;
                  Type_Sel_7     <=  3'b000;
                  Bypass_Sel_0   <=  3'b000;
                  Bypass_Sel_1   <=  3'b000;
                  Bypass_Sel_2   <=  3'b000;
                  Bypass_Sel_3   <=  3'b000;
                  Bypass_Sel_4   <=  3'b000;
                  Bypass_Sel_5   <=  3'b000;
                  Bypass_Sel_6   <=  3'b000;
                  Bypass_Sel_7   <=  3'b000;
                  DeShuf_Ctrl_0  <=  3'b000;
                  DeShuf_Ctrl_1  <=  3'b000;
                  DeShuf_Ctrl_2  <=  3'b000;
                  DeShuf_Ctrl_3  <=  3'b000;
                  DeShuf_Ctrl_4  <=  3'b000;
                  DeShuf_Ctrl_5  <=  3'b000;
                  DeShuf_Ctrl_6  <=  3'b000;
                  DeShuf_Ctrl_7  <=  3'b000;
                  Bypass_EN_0    <=  1'b0;
                  Bypass_EN_1    <=  1'b0;
                  Bypass_EN_2    <=  1'b0;
                  Bypass_EN_3    <=  1'b0;
                  Bypass_EN_4    <=  1'b0;
                  Bypass_EN_5    <=  1'b0;
                  Bypass_EN_6    <=  1'b0;
                  Bypass_EN_7    <=  1'b0;
                  Hold_Ctrl_0    <=  1'b0;
                  Hold_Ctrl_1    <=  1'b0;
                  Hold_Ctrl_2    <=  1'b0;
                  Hold_Ctrl_3    <=  1'b0;
                  Hold_Ctrl_4    <=  1'b0;
                  Hold_Ctrl_5    <=  1'b0;
                  Hold_Ctrl_6    <=  1'b0;
                  Hold_Ctrl_7    <=  1'b0;
                  DFF_Ctrl_0     <=  1'b0;
                  DFF_Ctrl_1     <=  1'b0;
                  DFF_Ctrl_2     <=  1'b0;
                  DFF_Ctrl_3     <=  1'b0;
                  DFF_Ctrl_4     <=  1'b0;
                  DFF_Ctrl_5     <=  1'b0;
                  DFF_Ctrl_6     <=  1'b0;
                  DFF_Ctrl_7     <=  1'b0;
                  hold_seg_0     <=  1'b0;
                  hold_seg_1     <=  1'b0;
                  hold_seg_2     <=  1'b0;
                  hold_seg_3     <=  1'b0;
                  hold_seg_4     <=  1'b0;
                  hold_seg_5     <=  1'b0;
                  hold_seg_6     <=  1'b0;
                  hold_seg_7     <=  1'b0;
                  in_ctrl_all_cb <=  1'b0;
                  hold_all_out   <=  1'b0;
                  in_ctrl_all_out<=  1'b1;
                  counter_en     <=  1'b1;
                  currentstate   <= state_15;
                end
              state_15:
                begin
                  hold_all_in    <=  1'b0;
                  hold_buf_2     <=  1'b1;
                  hold_buf_1     <=  1'b1;
                  hold_buf_0     <=  1'b1;
                  in_ctrl_buf_2  <=  1'b0;
                  in_ctrl_buf_1  <=  1'b0;
                  in_ctrl_buf_0  <=  1'b0;
                  pos_hold_ctrl  <=  1'b0;
                  Shuf_Ctrl_0    <=  3'b000;
                  Shuf_Ctrl_1    <=  3'b000;
                  Shuf_Ctrl_2    <=  3'b000;
                  Shuf_Ctrl_3    <=  3'b000;
                  Shuf_Ctrl_4    <=  3'b000;
                  Shuf_Ctrl_5    <=  3'b000;
                  Shuf_Ctrl_6    <=  3'b000;
                  Shuf_Ctrl_7    <=  3'b000;
                  Type_Sel_0     <=  3'b000;
                  Type_Sel_1     <=  3'b000;
                  Type_Sel_2     <=  3'b000;
                  Type_Sel_3     <=  3'b000;
                  Type_Sel_4     <=  3'b000;
                  Type_Sel_5     <=  3'b000;
                  Type_Sel_6     <=  3'b000;
                  Type_Sel_7     <=  3'b000;
                  Bypass_Sel_0   <=  3'b000;
                  Bypass_Sel_1   <=  3'b000;
                  Bypass_Sel_2   <=  3'b000;
                  Bypass_Sel_3   <=  3'b000;
                  Bypass_Sel_4   <=  3'b000;
                  Bypass_Sel_5   <=  3'b000;
                  Bypass_Sel_6   <=  3'b000;
                  Bypass_Sel_7   <=  3'b000;
                  DeShuf_Ctrl_0  <=  3'b000;
                  DeShuf_Ctrl_1  <=  3'b000;
                  DeShuf_Ctrl_2  <=  3'b000;
                  DeShuf_Ctrl_3  <=  3'b000;
                  DeShuf_Ctrl_4  <=  3'b000;
                  DeShuf_Ctrl_5  <=  3'b000;
                  DeShuf_Ctrl_6  <=  3'b000;
                  DeShuf_Ctrl_7  <=  3'b000;
                  Bypass_EN_0    <=  1'b0;
                  Bypass_EN_1    <=  1'b0;
                  Bypass_EN_2    <=  1'b0;
                  Bypass_EN_3    <=  1'b0;
                  Bypass_EN_4    <=  1'b0;
                  Bypass_EN_5    <=  1'b0;
                  Bypass_EN_6    <=  1'b0;
                  Bypass_EN_7    <=  1'b0;
                  Hold_Ctrl_0    <=  1'b0;
                  Hold_Ctrl_1    <=  1'b0;
                  Hold_Ctrl_2    <=  1'b0;
                  Hold_Ctrl_3    <=  1'b0;
                  Hold_Ctrl_4    <=  1'b0;
                  Hold_Ctrl_5    <=  1'b0;
                  Hold_Ctrl_6    <=  1'b0;
                  Hold_Ctrl_7    <=  1'b0;
                  DFF_Ctrl_0     <=  1'b0;
                  DFF_Ctrl_1     <=  1'b0;
                  DFF_Ctrl_2     <=  1'b0;
                  DFF_Ctrl_3     <=  1'b0;
                  DFF_Ctrl_4     <=  1'b0;
                  DFF_Ctrl_5     <=  1'b0;
                  DFF_Ctrl_6     <=  1'b0;
                  DFF_Ctrl_7     <=  1'b0;
                  hold_seg_0     <=  1'b0;
                  hold_seg_1     <=  1'b0;
                  hold_seg_2     <=  1'b0;
                  hold_seg_3     <=  1'b0;
                  hold_seg_4     <=  1'b0;
                  hold_seg_5     <=  1'b0;
                  hold_seg_6     <=  1'b0;
                  hold_seg_7     <=  1'b0;
                  in_ctrl_all_cb <=  1'b0;
                  hold_all_out   <=  1'b0;
                  in_ctrl_all_out<=  1'b1;
                  counter_en     <=  1'b0;
                  currentstate   <= state_16;
                end
              state_16:
                begin
                  hold_all_in    <=  1'b0;
                  hold_buf_2     <=  1'b1;
                  hold_buf_1     <=  1'b1;
                  hold_buf_0     <=  1'b1;
                  in_ctrl_buf_2  <=  1'b0;
                  in_ctrl_buf_1  <=  1'b0;
                  in_ctrl_buf_0  <=  1'b0;
                  pos_hold_ctrl  <=  1'b0;
                  Shuf_Ctrl_0    <=  3'b000;
                  Shuf_Ctrl_1    <=  3'b000;
                  Shuf_Ctrl_2    <=  3'b000;
                  Shuf_Ctrl_3    <=  3'b000;
                  Shuf_Ctrl_4    <=  3'b000;
                  Shuf_Ctrl_5    <=  3'b000;
                  Shuf_Ctrl_6    <=  3'b000;
                  Shuf_Ctrl_7    <=  3'b000;
                  Type_Sel_0     <=  3'b000;
                  Type_Sel_1     <=  3'b000;
                  Type_Sel_2     <=  3'b000;
                  Type_Sel_3     <=  3'b000;
                  Type_Sel_4     <=  3'b000;
                  Type_Sel_5     <=  3'b000;
                  Type_Sel_6     <=  3'b000;
                  Type_Sel_7     <=  3'b000;
                  Bypass_Sel_0   <=  3'b000;
                  Bypass_Sel_1   <=  3'b000;
                  Bypass_Sel_2   <=  3'b000;
                  Bypass_Sel_3   <=  3'b000;
                  Bypass_Sel_4   <=  3'b000;
                  Bypass_Sel_5   <=  3'b000;
                  Bypass_Sel_6   <=  3'b000;
                  Bypass_Sel_7   <=  3'b000;
                  DeShuf_Ctrl_0  <=  3'b000;
                  DeShuf_Ctrl_1  <=  3'b000;
                  DeShuf_Ctrl_2  <=  3'b000;
                  DeShuf_Ctrl_3  <=  3'b000;
                  DeShuf_Ctrl_4  <=  3'b000;
                  DeShuf_Ctrl_5  <=  3'b000;
                  DeShuf_Ctrl_6  <=  3'b000;
                  DeShuf_Ctrl_7  <=  3'b000;
                  Bypass_EN_0    <=  1'b0;
                  Bypass_EN_1    <=  1'b0;
                  Bypass_EN_2    <=  1'b0;
                  Bypass_EN_3    <=  1'b0;
                  Bypass_EN_4    <=  1'b0;
                  Bypass_EN_5    <=  1'b0;
                  Bypass_EN_6    <=  1'b0;
                  Bypass_EN_7    <=  1'b0;
                  Hold_Ctrl_0    <=  1'b0;
                  Hold_Ctrl_1    <=  1'b0;
                  Hold_Ctrl_2    <=  1'b0;
                  Hold_Ctrl_3    <=  1'b0;
                  Hold_Ctrl_4    <=  1'b0;
                  Hold_Ctrl_5    <=  1'b0;
                  Hold_Ctrl_6    <=  1'b0;
                  Hold_Ctrl_7    <=  1'b0;
                  DFF_Ctrl_0     <=  1'b0;
                  DFF_Ctrl_1     <=  1'b0;
                  DFF_Ctrl_2     <=  1'b0;
                  DFF_Ctrl_3     <=  1'b0;
                  DFF_Ctrl_4     <=  1'b0;
                  DFF_Ctrl_5     <=  1'b0;
                  DFF_Ctrl_6     <=  1'b0;
                  DFF_Ctrl_7     <=  1'b0;
                  hold_seg_0     <=  1'b0;
                  hold_seg_1     <=  1'b0;
                  hold_seg_2     <=  1'b0;
                  hold_seg_3     <=  1'b0;
                  hold_seg_4     <=  1'b0;
                  hold_seg_5     <=  1'b0;
                  hold_seg_6     <=  1'b0;
                  hold_seg_7     <=  1'b0;
                  in_ctrl_all_cb <=  1'b0;
                  hold_all_out   <=  1'b0;
                  in_ctrl_all_out<=  1'b1;
                  counter_en     <=  1'b0;
                  currentstate   <= state_17;
                end
              state_17:
                begin
                  hold_all_in    <=  1'b0;
                  hold_buf_2     <=  1'b1;
                  hold_buf_1     <=  1'b1;
                  hold_buf_0     <=  1'b1;
                  in_ctrl_buf_2  <=  1'b0;
                  in_ctrl_buf_1  <=  1'b0;
                  in_ctrl_buf_0  <=  1'b0;
                  pos_hold_ctrl  <=  1'b0;
                  Shuf_Ctrl_0    <=  3'b000;
                  Shuf_Ctrl_1    <=  3'b000;
                  Shuf_Ctrl_2    <=  3'b000;
                  Shuf_Ctrl_3    <=  3'b000;
                  Shuf_Ctrl_4    <=  3'b000;
                  Shuf_Ctrl_5    <=  3'b000;
                  Shuf_Ctrl_6    <=  3'b000;
                  Shuf_Ctrl_7    <=  3'b000;
                  Type_Sel_0     <=  3'b000;
                  Type_Sel_1     <=  3'b000;
                  Type_Sel_2     <=  3'b000;
                  Type_Sel_3     <=  3'b000;
                  Type_Sel_4     <=  3'b000;
                  Type_Sel_5     <=  3'b000;
                  Type_Sel_6     <=  3'b000;
                  Type_Sel_7     <=  3'b000;
                  Bypass_Sel_0   <=  3'b000;
                  Bypass_Sel_1   <=  3'b000;
                  Bypass_Sel_2   <=  3'b000;
                  Bypass_Sel_3   <=  3'b000;
                  Bypass_Sel_4   <=  3'b000;
                  Bypass_Sel_5   <=  3'b000;
                  Bypass_Sel_6   <=  3'b000;
                  Bypass_Sel_7   <=  3'b000;
                  DeShuf_Ctrl_0  <=  3'b000;
                  DeShuf_Ctrl_1  <=  3'b000;
                  DeShuf_Ctrl_2  <=  3'b000;
                  DeShuf_Ctrl_3  <=  3'b000;
                  DeShuf_Ctrl_4  <=  3'b000;
                  DeShuf_Ctrl_5  <=  3'b000;
                  DeShuf_Ctrl_6  <=  3'b000;
                  DeShuf_Ctrl_7  <=  3'b000;
                  Bypass_EN_0    <=  1'b0;
                  Bypass_EN_1    <=  1'b0;
                  Bypass_EN_2    <=  1'b0;
                  Bypass_EN_3    <=  1'b0;
                  Bypass_EN_4    <=  1'b0;
                  Bypass_EN_5    <=  1'b0;
                  Bypass_EN_6    <=  1'b0;
                  Bypass_EN_7    <=  1'b0;
                  Hold_Ctrl_0    <=  1'b0;
                  Hold_Ctrl_1    <=  1'b0;
                  Hold_Ctrl_2    <=  1'b0;
                  Hold_Ctrl_3    <=  1'b0;
                  Hold_Ctrl_4    <=  1'b0;
                  Hold_Ctrl_5    <=  1'b0;
                  Hold_Ctrl_6    <=  1'b0;
                  Hold_Ctrl_7    <=  1'b0;
                  DFF_Ctrl_0     <=  1'b0;
                  DFF_Ctrl_1     <=  1'b0;
                  DFF_Ctrl_2     <=  1'b0;
                  DFF_Ctrl_3     <=  1'b0;
                  DFF_Ctrl_4     <=  1'b0;
                  DFF_Ctrl_5     <=  1'b0;
                  DFF_Ctrl_6     <=  1'b0;
                  DFF_Ctrl_7     <=  1'b0;
                  hold_seg_0     <=  1'b0;
                  hold_seg_1     <=  1'b0;
                  hold_seg_2     <=  1'b0;
                  hold_seg_3     <=  1'b0;
                  hold_seg_4     <=  1'b0;
                  hold_seg_5     <=  1'b0;
                  hold_seg_6     <=  1'b0;
                  hold_seg_7     <=  1'b0;
                  in_ctrl_all_cb <=  1'b0;
                  hold_all_out   <=  1'b0;
                  in_ctrl_all_out<=  1'b1;
                  counter_en     <=  1'b0;
                  currentstate   <= state_18;
                end
              state_18:
                begin
                  hold_all_in    <=  1'b0;
                  hold_buf_2     <=  1'b1;
                  hold_buf_1     <=  1'b1;
                  hold_buf_0     <=  1'b1;
                  in_ctrl_buf_2  <=  1'b0;
                  in_ctrl_buf_1  <=  1'b0;
                  in_ctrl_buf_0  <=  1'b0;
                  pos_hold_ctrl  <=  1'b0;
                  Shuf_Ctrl_0    <=  3'b000;
                  Shuf_Ctrl_1    <=  3'b000;
                  Shuf_Ctrl_2    <=  3'b000;
                  Shuf_Ctrl_3    <=  3'b000;
                  Shuf_Ctrl_4    <=  3'b000;
                  Shuf_Ctrl_5    <=  3'b000;
                  Shuf_Ctrl_6    <=  3'b000;
                  Shuf_Ctrl_7    <=  3'b000;
                  Type_Sel_0     <=  3'b000;
                  Type_Sel_1     <=  3'b000;
                  Type_Sel_2     <=  3'b000;
                  Type_Sel_3     <=  3'b000;
                  Type_Sel_4     <=  3'b000;
                  Type_Sel_5     <=  3'b000;
                  Type_Sel_6     <=  3'b000;
                  Type_Sel_7     <=  3'b000;
                  Bypass_Sel_0   <=  3'b000;
                  Bypass_Sel_1   <=  3'b000;
                  Bypass_Sel_2   <=  3'b000;
                  Bypass_Sel_3   <=  3'b000;
                  Bypass_Sel_4   <=  3'b000;
                  Bypass_Sel_5   <=  3'b000;
                  Bypass_Sel_6   <=  3'b000;
                  Bypass_Sel_7   <=  3'b000;
                  DeShuf_Ctrl_0  <=  3'b000;
                  DeShuf_Ctrl_1  <=  3'b000;
                  DeShuf_Ctrl_2  <=  3'b000;
                  DeShuf_Ctrl_3  <=  3'b000;
                  DeShuf_Ctrl_4  <=  3'b000;
                  DeShuf_Ctrl_5  <=  3'b000;
                  DeShuf_Ctrl_6  <=  3'b000;
                  DeShuf_Ctrl_7  <=  3'b000;
                  Bypass_EN_0    <=  1'b0;
                  Bypass_EN_1    <=  1'b0;
                  Bypass_EN_2    <=  1'b0;
                  Bypass_EN_3    <=  1'b0;
                  Bypass_EN_4    <=  1'b0;
                  Bypass_EN_5    <=  1'b0;
                  Bypass_EN_6    <=  1'b0;
                  Bypass_EN_7    <=  1'b0;
                  Hold_Ctrl_0    <=  1'b0;
                  Hold_Ctrl_1    <=  1'b0;
                  Hold_Ctrl_2    <=  1'b0;
                  Hold_Ctrl_3    <=  1'b0;
                  Hold_Ctrl_4    <=  1'b0;
                  Hold_Ctrl_5    <=  1'b0;
                  Hold_Ctrl_6    <=  1'b0;
                  Hold_Ctrl_7    <=  1'b0;
                  DFF_Ctrl_0     <=  1'b0;
                  DFF_Ctrl_1     <=  1'b0;
                  DFF_Ctrl_2     <=  1'b0;
                  DFF_Ctrl_3     <=  1'b0;
                  DFF_Ctrl_4     <=  1'b0;
                  DFF_Ctrl_5     <=  1'b0;
                  DFF_Ctrl_6     <=  1'b0;
                  DFF_Ctrl_7     <=  1'b0;
                  hold_seg_0     <=  1'b0;
                  hold_seg_1     <=  1'b0;
                  hold_seg_2     <=  1'b0;
                  hold_seg_3     <=  1'b0;
                  hold_seg_4     <=  1'b0;
                  hold_seg_5     <=  1'b0;
                  hold_seg_6     <=  1'b0;
                  hold_seg_7     <=  1'b0;
                  in_ctrl_all_cb <=  1'b0;
                  hold_all_out   <=  1'b0;
                  in_ctrl_all_out<=  1'b1;
                  counter_en     <=  1'b0;
                  currentstate   <= state_19;
                end
              state_19:
                begin
                  hold_all_in    <=  1'b0;
                  hold_buf_2     <=  1'b1;
                  hold_buf_1     <=  1'b1;
                  hold_buf_0     <=  1'b1;
                  in_ctrl_buf_2  <=  1'b0;
                  in_ctrl_buf_1  <=  1'b0;
                  in_ctrl_buf_0  <=  1'b0;
                  pos_hold_ctrl  <=  1'b0;
                  Shuf_Ctrl_0    <=  3'b000;
                  Shuf_Ctrl_1    <=  3'b000;
                  Shuf_Ctrl_2    <=  3'b000;
                  Shuf_Ctrl_3    <=  3'b000;
                  Shuf_Ctrl_4    <=  3'b000;
                  Shuf_Ctrl_5    <=  3'b000;
                  Shuf_Ctrl_6    <=  3'b000;
                  Shuf_Ctrl_7    <=  3'b000;
                  Type_Sel_0     <=  3'b000;
                  Type_Sel_1     <=  3'b000;
                  Type_Sel_2     <=  3'b000;
                  Type_Sel_3     <=  3'b000;
                  Type_Sel_4     <=  3'b000;
                  Type_Sel_5     <=  3'b000;
                  Type_Sel_6     <=  3'b000;
                  Type_Sel_7     <=  3'b000;
                  Bypass_Sel_0   <=  3'b000;
                  Bypass_Sel_1   <=  3'b000;
                  Bypass_Sel_2   <=  3'b000;
                  Bypass_Sel_3   <=  3'b000;
                  Bypass_Sel_4   <=  3'b000;
                  Bypass_Sel_5   <=  3'b000;
                  Bypass_Sel_6   <=  3'b000;
                  Bypass_Sel_7   <=  3'b000;
                  DeShuf_Ctrl_0  <=  3'b000;
                  DeShuf_Ctrl_1  <=  3'b000;
                  DeShuf_Ctrl_2  <=  3'b000;
                  DeShuf_Ctrl_3  <=  3'b000;
                  DeShuf_Ctrl_4  <=  3'b000;
                  DeShuf_Ctrl_5  <=  3'b000;
                  DeShuf_Ctrl_6  <=  3'b000;
                  DeShuf_Ctrl_7  <=  3'b000;
                  Bypass_EN_0    <=  1'b0;
                  Bypass_EN_1    <=  1'b0;
                  Bypass_EN_2    <=  1'b0;
                  Bypass_EN_3    <=  1'b0;
                  Bypass_EN_4    <=  1'b0;
                  Bypass_EN_5    <=  1'b0;
                  Bypass_EN_6    <=  1'b0;
                  Bypass_EN_7    <=  1'b0;
                  Hold_Ctrl_0    <=  1'b0;
                  Hold_Ctrl_1    <=  1'b0;
                  Hold_Ctrl_2    <=  1'b0;
                  Hold_Ctrl_3    <=  1'b0;
                  Hold_Ctrl_4    <=  1'b0;
                  Hold_Ctrl_5    <=  1'b0;
                  Hold_Ctrl_6    <=  1'b0;
                  Hold_Ctrl_7    <=  1'b0;
                  DFF_Ctrl_0     <=  1'b0;
                  DFF_Ctrl_1     <=  1'b0;
                  DFF_Ctrl_2     <=  1'b0;
                  DFF_Ctrl_3     <=  1'b0;
                  DFF_Ctrl_4     <=  1'b0;
                  DFF_Ctrl_5     <=  1'b0;
                  DFF_Ctrl_6     <=  1'b0;
                  DFF_Ctrl_7     <=  1'b0;
                  hold_seg_0     <=  1'b0;
                  hold_seg_1     <=  1'b0;
                  hold_seg_2     <=  1'b0;
                  hold_seg_3     <=  1'b0;
                  hold_seg_4     <=  1'b0;
                  hold_seg_5     <=  1'b0;
                  hold_seg_6     <=  1'b0;
                  hold_seg_7     <=  1'b0;
                  in_ctrl_all_cb <=  1'b0;
                  hold_all_out   <=  1'b0;
                  in_ctrl_all_out<=  1'b1;
                  counter_en     <=  1'b0;
                  currentstate   <= state_20;
                end
              state_20:
                begin
                  hold_all_in    <=  1'b0;
                  hold_buf_2     <=  1'b1;
                  hold_buf_1     <=  1'b1;
                  hold_buf_0     <=  1'b1;
                  in_ctrl_buf_2  <=  1'b0;
                  in_ctrl_buf_1  <=  1'b0;
                  in_ctrl_buf_0  <=  1'b0;
                  pos_hold_ctrl  <=  1'b0;
                  Shuf_Ctrl_0    <=  3'b000;
                  Shuf_Ctrl_1    <=  3'b000;
                  Shuf_Ctrl_2    <=  3'b000;
                  Shuf_Ctrl_3    <=  3'b000;
                  Shuf_Ctrl_4    <=  3'b000;
                  Shuf_Ctrl_5    <=  3'b000;
                  Shuf_Ctrl_6    <=  3'b000;
                  Shuf_Ctrl_7    <=  3'b000;
                  Type_Sel_0     <=  3'b000;
                  Type_Sel_1     <=  3'b000;
                  Type_Sel_2     <=  3'b000;
                  Type_Sel_3     <=  3'b000;
                  Type_Sel_4     <=  3'b000;
                  Type_Sel_5     <=  3'b000;
                  Type_Sel_6     <=  3'b000;
                  Type_Sel_7     <=  3'b000;
                  Bypass_Sel_0   <=  3'b000;
                  Bypass_Sel_1   <=  3'b000;
                  Bypass_Sel_2   <=  3'b000;
                  Bypass_Sel_3   <=  3'b000;
                  Bypass_Sel_4   <=  3'b000;
                  Bypass_Sel_5   <=  3'b000;
                  Bypass_Sel_6   <=  3'b000;
                  Bypass_Sel_7   <=  3'b000;
                  DeShuf_Ctrl_0  <=  3'b000;
                  DeShuf_Ctrl_1  <=  3'b000;
                  DeShuf_Ctrl_2  <=  3'b000;
                  DeShuf_Ctrl_3  <=  3'b000;
                  DeShuf_Ctrl_4  <=  3'b000;
                  DeShuf_Ctrl_5  <=  3'b000;
                  DeShuf_Ctrl_6  <=  3'b000;
                  DeShuf_Ctrl_7  <=  3'b000;
                  Bypass_EN_0    <=  1'b0;
                  Bypass_EN_1    <=  1'b0;
                  Bypass_EN_2    <=  1'b0;
                  Bypass_EN_3    <=  1'b0;
                  Bypass_EN_4    <=  1'b0;
                  Bypass_EN_5    <=  1'b0;
                  Bypass_EN_6    <=  1'b0;
                  Bypass_EN_7    <=  1'b0;
                  Hold_Ctrl_0    <=  1'b0;
                  Hold_Ctrl_1    <=  1'b0;
                  Hold_Ctrl_2    <=  1'b0;
                  Hold_Ctrl_3    <=  1'b0;
                  Hold_Ctrl_4    <=  1'b0;
                  Hold_Ctrl_5    <=  1'b0;
                  Hold_Ctrl_6    <=  1'b0;
                  Hold_Ctrl_7    <=  1'b0;
                  DFF_Ctrl_0     <=  1'b0;
                  DFF_Ctrl_1     <=  1'b0;
                  DFF_Ctrl_2     <=  1'b0;
                  DFF_Ctrl_3     <=  1'b0;
                  DFF_Ctrl_4     <=  1'b0;
                  DFF_Ctrl_5     <=  1'b0;
                  DFF_Ctrl_6     <=  1'b0;
                  DFF_Ctrl_7     <=  1'b0;
                  hold_seg_0     <=  1'b0;
                  hold_seg_1     <=  1'b0;
                  hold_seg_2     <=  1'b0;
                  hold_seg_3     <=  1'b0;
                  hold_seg_4     <=  1'b0;
                  hold_seg_5     <=  1'b0;
                  hold_seg_6     <=  1'b0;
                  hold_seg_7     <=  1'b0;
                  in_ctrl_all_cb <=  1'b0;
                  hold_all_out   <=  1'b0;
                  in_ctrl_all_out<=  1'b1;
                  counter_en     <=  1'b0;
                  currentstate   <= state_21;
                end
              state_21:
                begin
                  hold_all_in    <=  1'b0;
                  hold_buf_2     <=  1'b1;
                  hold_buf_1     <=  1'b1;
                  hold_buf_0     <=  1'b1;
                  in_ctrl_buf_2  <=  1'b0;
                  in_ctrl_buf_1  <=  1'b0;
                  in_ctrl_buf_0  <=  1'b0;
                  pos_hold_ctrl  <=  1'b0;
                  Shuf_Ctrl_0    <=  3'b000;
                  Shuf_Ctrl_1    <=  3'b000;
                  Shuf_Ctrl_2    <=  3'b000;
                  Shuf_Ctrl_3    <=  3'b000;
                  Shuf_Ctrl_4    <=  3'b000;
                  Shuf_Ctrl_5    <=  3'b000;
                  Shuf_Ctrl_6    <=  3'b000;
                  Shuf_Ctrl_7    <=  3'b000;
                  Type_Sel_0     <=  3'b000;
                  Type_Sel_1     <=  3'b000;
                  Type_Sel_2     <=  3'b000;
                  Type_Sel_3     <=  3'b000;
                  Type_Sel_4     <=  3'b000;
                  Type_Sel_5     <=  3'b000;
                  Type_Sel_6     <=  3'b000;
                  Type_Sel_7     <=  3'b000;
                  Bypass_Sel_0   <=  3'b000;
                  Bypass_Sel_1   <=  3'b000;
                  Bypass_Sel_2   <=  3'b000;
                  Bypass_Sel_3   <=  3'b000;
                  Bypass_Sel_4   <=  3'b000;
                  Bypass_Sel_5   <=  3'b000;
                  Bypass_Sel_6   <=  3'b000;
                  Bypass_Sel_7   <=  3'b000;
                  DeShuf_Ctrl_0  <=  3'b000;
                  DeShuf_Ctrl_1  <=  3'b000;
                  DeShuf_Ctrl_2  <=  3'b000;
                  DeShuf_Ctrl_3  <=  3'b000;
                  DeShuf_Ctrl_4  <=  3'b000;
                  DeShuf_Ctrl_5  <=  3'b000;
                  DeShuf_Ctrl_6  <=  3'b000;
                  DeShuf_Ctrl_7  <=  3'b000;
                  Bypass_EN_0    <=  1'b0;
                  Bypass_EN_1    <=  1'b0;
                  Bypass_EN_2    <=  1'b0;
                  Bypass_EN_3    <=  1'b0;
                  Bypass_EN_4    <=  1'b0;
                  Bypass_EN_5    <=  1'b0;
                  Bypass_EN_6    <=  1'b0;
                  Bypass_EN_7    <=  1'b0;
                  Hold_Ctrl_0    <=  1'b0;
                  Hold_Ctrl_1    <=  1'b0;
                  Hold_Ctrl_2    <=  1'b0;
                  Hold_Ctrl_3    <=  1'b0;
                  Hold_Ctrl_4    <=  1'b0;
                  Hold_Ctrl_5    <=  1'b0;
                  Hold_Ctrl_6    <=  1'b0;
                  Hold_Ctrl_7    <=  1'b0;
                  DFF_Ctrl_0     <=  1'b0;
                  DFF_Ctrl_1     <=  1'b0;
                  DFF_Ctrl_2     <=  1'b0;
                  DFF_Ctrl_3     <=  1'b0;
                  DFF_Ctrl_4     <=  1'b0;
                  DFF_Ctrl_5     <=  1'b0;
                  DFF_Ctrl_6     <=  1'b0;
                  DFF_Ctrl_7     <=  1'b0;
                  hold_seg_0     <=  1'b0;
                  hold_seg_1     <=  1'b0;
                  hold_seg_2     <=  1'b0;
                  hold_seg_3     <=  1'b0;
                  hold_seg_4     <=  1'b0;
                  hold_seg_5     <=  1'b0;
                  hold_seg_6     <=  1'b0;
                  hold_seg_7     <=  1'b0;
                  in_ctrl_all_cb <=  1'b0;
                  hold_all_out   <=  1'b0;
                  in_ctrl_all_out<=  1'b0;
                  counter_en     <=  1'b0;
                  currentstate   <= state_22;
                end
              state_22:
                begin
                  hold_all_in    <=  1'b0;
                  hold_buf_2     <=  1'b1;
                  hold_buf_1     <=  1'b1;
                  hold_buf_0     <=  1'b1;
                  in_ctrl_buf_2  <=  1'b0;
                  in_ctrl_buf_1  <=  1'b0;
                  in_ctrl_buf_0  <=  1'b0;
                  pos_hold_ctrl  <=  1'b0;
                  Shuf_Ctrl_0    <=  3'b000;
                  Shuf_Ctrl_1    <=  3'b000;
                  Shuf_Ctrl_2    <=  3'b000;
                  Shuf_Ctrl_3    <=  3'b000;
                  Shuf_Ctrl_4    <=  3'b000;
                  Shuf_Ctrl_5    <=  3'b000;
                  Shuf_Ctrl_6    <=  3'b000;
                  Shuf_Ctrl_7    <=  3'b000;
                  Type_Sel_0     <=  3'b000;
                  Type_Sel_1     <=  3'b000;
                  Type_Sel_2     <=  3'b000;
                  Type_Sel_3     <=  3'b000;
                  Type_Sel_4     <=  3'b000;
                  Type_Sel_5     <=  3'b000;
                  Type_Sel_6     <=  3'b000;
                  Type_Sel_7     <=  3'b000;
                  Bypass_Sel_0   <=  3'b000;
                  Bypass_Sel_1   <=  3'b000;
                  Bypass_Sel_2   <=  3'b000;
                  Bypass_Sel_3   <=  3'b000;
                  Bypass_Sel_4   <=  3'b000;
                  Bypass_Sel_5   <=  3'b000;
                  Bypass_Sel_6   <=  3'b000;
                  Bypass_Sel_7   <=  3'b000;
                  DeShuf_Ctrl_0  <=  3'b000;
                  DeShuf_Ctrl_1  <=  3'b000;
                  DeShuf_Ctrl_2  <=  3'b000;
                  DeShuf_Ctrl_3  <=  3'b000;
                  DeShuf_Ctrl_4  <=  3'b000;
                  DeShuf_Ctrl_5  <=  3'b000;
                  DeShuf_Ctrl_6  <=  3'b000;
                  DeShuf_Ctrl_7  <=  3'b000;
                  Bypass_EN_0    <=  1'b0;
                  Bypass_EN_1    <=  1'b0;
                  Bypass_EN_2    <=  1'b0;
                  Bypass_EN_3    <=  1'b0;
                  Bypass_EN_4    <=  1'b0;
                  Bypass_EN_5    <=  1'b0;
                  Bypass_EN_6    <=  1'b0;
                  Bypass_EN_7    <=  1'b0;
                  Hold_Ctrl_0    <=  1'b0;
                  Hold_Ctrl_1    <=  1'b0;
                  Hold_Ctrl_2    <=  1'b0;
                  Hold_Ctrl_3    <=  1'b0;
                  Hold_Ctrl_4    <=  1'b0;
                  Hold_Ctrl_5    <=  1'b0;
                  Hold_Ctrl_6    <=  1'b0;
                  Hold_Ctrl_7    <=  1'b0;
                  DFF_Ctrl_0     <=  1'b0;
                  DFF_Ctrl_1     <=  1'b0;
                  DFF_Ctrl_2     <=  1'b0;
                  DFF_Ctrl_3     <=  1'b0;
                  DFF_Ctrl_4     <=  1'b0;
                  DFF_Ctrl_5     <=  1'b0;
                  DFF_Ctrl_6     <=  1'b0;
                  DFF_Ctrl_7     <=  1'b0;
                  hold_seg_0     <=  1'b1;
                  hold_seg_1     <=  1'b1;
                  hold_seg_2     <=  1'b1;
                  hold_seg_3     <=  1'b1;
                  hold_seg_4     <=  1'b1;
                  hold_seg_5     <=  1'b1;
                  hold_seg_6     <=  1'b1;
                  hold_seg_7     <=  1'b1;
                  in_ctrl_all_cb <=  1'b1;
                  hold_all_out   <=  1'b0;
                  in_ctrl_all_out<=  1'b0;
                  counter_en     <=  1'b0;
                  currentstate   <= state_0;
                end
          endcase
        end
    end
endmodule
