module complex_mult_twiddle_wn0_32b(
  A32,
  R32,
  );
  
   
  input  [31:0] A32;
  output [31:0] R32;


  assign R32 = A32;

endmodule
