LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY complex_subst_cla_32b IS
	PORT	(
				A32		:	IN	STD_LOGIC_VECTOR (31 DOWNTO 0);
				B32		:	IN	STD_LOGIC_VECTOR (31 DOWNTO 0);
				R32		:	OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
				C_OUT32	:	OUT STD_LOGIC_VECTOR (1 DOWNTO 0)
			);
END complex_subst_cla_32b;

ARCHITECTURE structural OF complex_subst_cla_32b IS
SIGNAL REAL_A32 : STD_LOGIC_VECTOR (15 DOWNTO 0);
SIGNAL REAL_B32 : STD_LOGIC_VECTOR (15 DOWNTO 0);
SIGNAL REAL_R32 : STD_LOGIC_VECTOR (15 DOWNTO 0);
SIGNAL IMAG_A32 : STD_LOGIC_VECTOR (15 DOWNTO 0);
SIGNAL IMAG_B32 : STD_LOGIC_VECTOR (15 DOWNTO 0);
SIGNAL IMAG_R32 : STD_LOGIC_VECTOR (15 DOWNTO 0);
COMPONENT subst_cla_16b IS
	PORT	(
				A16		:	IN	STD_LOGIC_VECTOR (15 DOWNTO 0);
				B16		:	IN	STD_LOGIC_VECTOR (15 DOWNTO 0);
				R16		:	OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
				C_OUT16	:	OUT STD_LOGIC
			);
END COMPONENT;
BEGIN
	REAL_A32			<= A32(31 DOWNTO 16);
	REAL_B32			<= B32(31 DOWNTO 16);
	IMAG_A32			<= A32(15 DOWNTO 0);
	IMAG_B32			<= B32(15 DOWNTO 0);
	R32(31 DOWNTO 16) 	<= REAL_R32;
	R32(15 DOWNTO 0)	<= IMAG_R32;
	ADDER_REAL	:
		subst_cla_16b
			PORT MAP 
				(
					A16		=>REAL_A32,
					B16		=>REAL_B32,
					R16		=>REAL_R32,
					C_OUT16 =>C_OUT32(1)
				);
	ADDER_IMAG	:
		subst_cla_16b
			PORT MAP 
				(
					A16		=>IMAG_A32,
					B16		=>IMAG_B32,
					R16		=>IMAG_R32,
					C_OUT16 =>C_OUT32(0)
				);
END structural;

