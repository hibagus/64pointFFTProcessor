LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;
USE ieee.std_logic_unsigned.all;

ENTITY master_control IS
	PORT	(
				clk		         : IN  STD_LOGIC;
			    rst		         : IN  STD_LOGIC;
				mastertrig		 : IN  STD_LOGIC;
                hold_all_in      : OUT STD_LOGIC;
                hold_buf_3       : OUT STD_LOGIC;
                hold_buf_2       : OUT STD_LOGIC;
                hold_buf_1       : OUT STD_LOGIC;
                in_ctrl_buf_3    : OUT STD_LOGIC;
                in_ctrl_buf_2    : OUT STD_LOGIC;
                in_ctrl_buf_1    : OUT STD_LOGIC;
                pos_hold_ctrl    : OUT STD_LOGIC;
                Shuf_Ctrl_1      : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
                Shuf_Ctrl_2      : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
                Shuf_Ctrl_3      : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
                Shuf_Ctrl_4      : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
                Shuf_Ctrl_5      : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
                Shuf_Ctrl_6      : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
                Shuf_Ctrl_7      : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
                Shuf_Ctrl_8      : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
                Type_Sel_1       : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
                Type_Sel_2       : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
                Type_Sel_3       : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
                Type_Sel_4       : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
                Type_Sel_5       : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
                Type_Sel_6       : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
                Type_Sel_7       : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
                Type_Sel_8       : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
                Bypass_Sel_0     : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
                Bypass_Sel_1     : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
                Bypass_Sel_2     : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
                Bypass_Sel_3     : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
                Bypass_Sel_4     : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
                Bypass_Sel_5     : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
                Bypass_Sel_6     : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
                Bypass_Sel_7     : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
                DeShuf_Ctrl_0    : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
                DeShuf_Ctrl_1    : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
                DeShuf_Ctrl_2    : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
                DeShuf_Ctrl_3    : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
                DeShuf_Ctrl_4    : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
                DeShuf_Ctrl_5    : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
                DeShuf_Ctrl_6    : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
                DeShuf_Ctrl_7    : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
                Bypass_EN_0      : OUT STD_LOGIC;
                Bypass_EN_1      : OUT STD_LOGIC;
                Bypass_EN_2      : OUT STD_LOGIC;
                Bypass_EN_3      : OUT STD_LOGIC;
                Bypass_EN_4      : OUT STD_LOGIC;
                Bypass_EN_5      : OUT STD_LOGIC;
                Bypass_EN_6      : OUT STD_LOGIC;
                Bypass_EN_7      : OUT STD_LOGIC;
                Hold_Ctrl_0      : OUT STD_LOGIC;
                Hold_Ctrl_1      : OUT STD_LOGIC;
                Hold_Ctrl_2      : OUT STD_LOGIC;
                Hold_Ctrl_3      : OUT STD_LOGIC;
                Hold_Ctrl_4      : OUT STD_LOGIC;
                Hold_Ctrl_5      : OUT STD_LOGIC;
                Hold_Ctrl_6      : OUT STD_LOGIC;
                Hold_Ctrl_7      : OUT STD_LOGIC;
                DFF_Ctrl_0       : OUT STD_LOGIC;
                DFF_Ctrl_1       : OUT STD_LOGIC;
                DFF_Ctrl_2       : OUT STD_LOGIC;
                DFF_Ctrl_3       : OUT STD_LOGIC;
                DFF_Ctrl_4       : OUT STD_LOGIC;
                DFF_Ctrl_5       : OUT STD_LOGIC;
                DFF_Ctrl_6       : OUT STD_LOGIC;
                DFF_Ctrl_7       : OUT STD_LOGIC;
                hold_seg_0       : OUT STD_LOGIC;
                hold_seg_1       : OUT STD_LOGIC;
                hold_seg_2       : OUT STD_LOGIC;
                hold_seg_3       : OUT STD_LOGIC;
                hold_seg_4       : OUT STD_LOGIC;
                hold_seg_5       : OUT STD_LOGIC;
                hold_seg_6       : OUT STD_LOGIC;
                hold_seg_7       : OUT STD_LOGIC;
                in_ctrl_all_cb   : OUT STD_LOGIC;
                hold_all_out     : OUT STD_LOGIC;
                in_ctrl_all_out  : OUT STD_LOGIC;
                counter_en       : OUT STD_LOGIC
			);
END master_control;

ARCHITECTURE behavioral OF master_control IS
TYPE FSMSTATE IS (
	state_0, state_1, state_2, state_3, state_4, state_5, state_6,  
	state_7, state_8, state_9, state_10, state_11, state_12, state_13, 
	state_14, state_15, state_16, state_17, state_18, state_19, state_20, 
	state_21, state_22
	);

SIGNAL currentstate	: FSMSTATE;
	BEGIN
	PROCESS(clk,rst,currentstate,mastertrig)
	BEGIN
		IF rst='1' THEN
			currentstate <= state_0;
		ELSE
			IF ((clk'EVENT) AND (clk='1'))  THEN
				CASE currentstate IS
                    WHEN state_0 		 =>
                        hold_all_in    <=  '0';
                        hold_buf_3     <=  '1';
                        hold_buf_2     <=  '1';
                        hold_buf_1     <=  '1';
                        in_ctrl_buf_3  <=  '0';
                        in_ctrl_buf_2  <=  '0';
                        in_ctrl_buf_1  <=  '0';
                        pos_hold_ctrl  <=  '0';
                        Shuf_Ctrl_1    <=  "000";
                        Shuf_Ctrl_2    <=  "000";
                        Shuf_Ctrl_3    <=  "000";
                        Shuf_Ctrl_4    <=  "000";
                        Shuf_Ctrl_5    <=  "000";
                        Shuf_Ctrl_6    <=  "000";
                        Shuf_Ctrl_7    <=  "000";
                        Shuf_Ctrl_8    <=  "000";
                        Type_Sel_1     <=  "000";
                        Type_Sel_2     <=  "000";
                        Type_Sel_3     <=  "000";
                        Type_Sel_4     <=  "000";
                        Type_Sel_5     <=  "000";
                        Type_Sel_6     <=  "000";
                        Type_Sel_7     <=  "000";
                        Type_Sel_8     <=  "000";
                        Bypass_Sel_0   <=  "000";
                        Bypass_Sel_1   <=  "000";
                        Bypass_Sel_2   <=  "000";
                        Bypass_Sel_3   <=  "000";
                        Bypass_Sel_4   <=  "000";
                        Bypass_Sel_5   <=  "000";
                        Bypass_Sel_6   <=  "000";
                        Bypass_Sel_7   <=  "000";
                        DeShuf_Ctrl_0  <=  "000";
                        DeShuf_Ctrl_1  <=  "000";
                        DeShuf_Ctrl_2  <=  "000";
                        DeShuf_Ctrl_3  <=  "000";
                        DeShuf_Ctrl_4  <=  "000";
                        DeShuf_Ctrl_5  <=  "000";
                        DeShuf_Ctrl_6  <=  "000";
                        DeShuf_Ctrl_7  <=  "000";
                        Bypass_EN_0    <=  '1';
                        Bypass_EN_1    <=  '1';
                        Bypass_EN_2    <=  '1';
                        Bypass_EN_3    <=  '1';
                        Bypass_EN_4    <=  '1';
                        Bypass_EN_5    <=  '1';
                        Bypass_EN_6    <=  '1';
                        Bypass_EN_7    <=  '1';
                        Hold_Ctrl_0    <=  '0';
                        Hold_Ctrl_1    <=  '0';
                        Hold_Ctrl_2    <=  '0';
                        Hold_Ctrl_3    <=  '0';
                        Hold_Ctrl_4    <=  '0';
                        Hold_Ctrl_5    <=  '0';
                        Hold_Ctrl_6    <=  '0';
                        Hold_Ctrl_7    <=  '0';
                        DFF_Ctrl_0     <=  '0';
                        DFF_Ctrl_1     <=  '0';
                        DFF_Ctrl_2     <=  '0';
                        DFF_Ctrl_3     <=  '0';
                        DFF_Ctrl_4     <=  '0';
                        DFF_Ctrl_5     <=  '0';
                        DFF_Ctrl_6     <=  '0';
                        DFF_Ctrl_7     <=  '0';
                        hold_seg_0     <=  '1';
                        hold_seg_1     <=  '1';
                        hold_seg_2     <=  '1';
                        hold_seg_3     <=  '1';
                        hold_seg_4     <=  '1';
                        hold_seg_5     <=  '1';
                        hold_seg_6     <=  '1';
                        hold_seg_7     <=  '1';
                        in_ctrl_all_cb <=  '1';
                        hold_all_out   <=  '0';
                        in_ctrl_all_out<=  '0';
                        counter_en     <=  '0';		
						IF mastertrig='1' THEN
							currentstate   <= state_1;
						ELSE
							currentstate   <= state_0;
						END IF;
                    WHEN state_1		 =>
                        hold_all_in    <=  '0';
                        hold_buf_3     <=  '1';
                        hold_buf_2     <=  '1';
                        hold_buf_1     <=  '1';
                        in_ctrl_buf_3  <=  '0';
                        in_ctrl_buf_2  <=  '0';
                        in_ctrl_buf_1  <=  '0';
                        pos_hold_ctrl  <=  '0';
                        Shuf_Ctrl_1    <=  "000";
                        Shuf_Ctrl_2    <=  "000";
                        Shuf_Ctrl_3    <=  "000";
                        Shuf_Ctrl_4    <=  "000";
                        Shuf_Ctrl_5    <=  "000";
                        Shuf_Ctrl_6    <=  "000";
                        Shuf_Ctrl_7    <=  "000";
                        Shuf_Ctrl_8    <=  "000";
                        Type_Sel_1     <=  "000";
                        Type_Sel_2     <=  "000";
                        Type_Sel_3     <=  "000";
                        Type_Sel_4     <=  "000";
                        Type_Sel_5     <=  "000";
                        Type_Sel_6     <=  "000";
                        Type_Sel_7     <=  "000";
                        Type_Sel_8     <=  "000";
                        Bypass_Sel_0   <=  "000";
                        Bypass_Sel_1   <=  "000";
                        Bypass_Sel_2   <=  "000";
                        Bypass_Sel_3   <=  "000";
                        Bypass_Sel_4   <=  "000";
                        Bypass_Sel_5   <=  "000";
                        Bypass_Sel_6   <=  "000";
                        Bypass_Sel_7   <=  "000";
                        DeShuf_Ctrl_0  <=  "000";
                        DeShuf_Ctrl_1  <=  "000";
                        DeShuf_Ctrl_2  <=  "000";
                        DeShuf_Ctrl_3  <=  "000";
                        DeShuf_Ctrl_4  <=  "000";
                        DeShuf_Ctrl_5  <=  "000";
                        DeShuf_Ctrl_6  <=  "000";
                        DeShuf_Ctrl_7  <=  "000";
                        Bypass_EN_0    <=  '1';
                        Bypass_EN_1    <=  '1';
                        Bypass_EN_2    <=  '1';
                        Bypass_EN_3    <=  '1';
                        Bypass_EN_4    <=  '1';
                        Bypass_EN_5    <=  '1';
                        Bypass_EN_6    <=  '1';
                        Bypass_EN_7    <=  '1';
                        Hold_Ctrl_0    <=  '0';
                        Hold_Ctrl_1    <=  '0';
                        Hold_Ctrl_2    <=  '0';
                        Hold_Ctrl_3    <=  '0';
                        Hold_Ctrl_4    <=  '0';
                        Hold_Ctrl_5    <=  '0';
                        Hold_Ctrl_6    <=  '0';
                        Hold_Ctrl_7    <=  '0';
                        DFF_Ctrl_0     <=  '0';
                        DFF_Ctrl_1     <=  '0';
                        DFF_Ctrl_2     <=  '0';
                        DFF_Ctrl_3     <=  '0';
                        DFF_Ctrl_4     <=  '0';
                        DFF_Ctrl_5     <=  '0';
                        DFF_Ctrl_6     <=  '0';
                        DFF_Ctrl_7     <=  '0';
                        hold_seg_0     <=  '0';
                        hold_seg_1     <=  '1';
                        hold_seg_2     <=  '1';
                        hold_seg_3     <=  '1';
                        hold_seg_4     <=  '1';
                        hold_seg_5     <=  '1';
                        hold_seg_6     <=  '1';
                        hold_seg_7     <=  '1';
                        in_ctrl_all_cb <=  '1';
                        hold_all_out   <=  '0';
                        in_ctrl_all_out<=  '0';
                        counter_en     <=  '0';
                        currentstate   <= state_2;					
                    WHEN state_2		 =>
                        hold_all_in    <=  '0';
                        hold_buf_3     <=  '1';
                        hold_buf_2     <=  '1';
                        hold_buf_1     <=  '1';
                        in_ctrl_buf_3  <=  '0';
                        in_ctrl_buf_2  <=  '0';
                        in_ctrl_buf_1  <=  '0';
                        pos_hold_ctrl  <=  '0';
                        Shuf_Ctrl_1    <=  "001";
                        Shuf_Ctrl_2    <=  "010";
                        Shuf_Ctrl_3    <=  "011";
                        Shuf_Ctrl_4    <=  "100";
                        Shuf_Ctrl_5    <=  "101";
                        Shuf_Ctrl_6    <=  "110";
                        Shuf_Ctrl_7    <=  "111";
                        Shuf_Ctrl_8    <=  "000";
                        Type_Sel_1     <=  "001";
                        Type_Sel_2     <=  "001";
                        Type_Sel_3     <=  "001";
                        Type_Sel_4     <=  "001";
                        Type_Sel_5     <=  "001";
                        Type_Sel_6     <=  "001";
                        Type_Sel_7     <=  "001";
                        Type_Sel_8     <=  "001";
                        Bypass_Sel_0   <=  "000";
                        Bypass_Sel_1   <=  "000";
                        Bypass_Sel_2   <=  "000";
                        Bypass_Sel_3   <=  "000";
                        Bypass_Sel_4   <=  "000";
                        Bypass_Sel_5   <=  "000";
                        Bypass_Sel_6   <=  "000";
                        Bypass_Sel_7   <=  "000";
                        DeShuf_Ctrl_0  <=  "000";
                        DeShuf_Ctrl_1  <=  "000";
                        DeShuf_Ctrl_2  <=  "001";
                        DeShuf_Ctrl_3  <=  "010";
                        DeShuf_Ctrl_4  <=  "011";
                        DeShuf_Ctrl_5  <=  "100";
                        DeShuf_Ctrl_6  <=  "101";
                        DeShuf_Ctrl_7  <=  "110";
                        Bypass_EN_0    <=  '1';
                        Bypass_EN_1    <=  '0';
                        Bypass_EN_2    <=  '0';
                        Bypass_EN_3    <=  '0';
                        Bypass_EN_4    <=  '0';
                        Bypass_EN_5    <=  '0';
                        Bypass_EN_6    <=  '0';
                        Bypass_EN_7    <=  '0';
                        Hold_Ctrl_0    <=  '0';
                        Hold_Ctrl_1    <=  '0';
                        Hold_Ctrl_2    <=  '0';
                        Hold_Ctrl_3    <=  '0';
                        Hold_Ctrl_4    <=  '0';
                        Hold_Ctrl_5    <=  '0';
                        Hold_Ctrl_6    <=  '0';
                        Hold_Ctrl_7    <=  '0';
                        DFF_Ctrl_0     <=  '0';
                        DFF_Ctrl_1     <=  '0';
                        DFF_Ctrl_2     <=  '0';
                        DFF_Ctrl_3     <=  '0';
                        DFF_Ctrl_4     <=  '0';
                        DFF_Ctrl_5     <=  '0';
                        DFF_Ctrl_6     <=  '0';
                        DFF_Ctrl_7     <=  '0';
                        hold_seg_0     <=  '1';
                        hold_seg_1     <=  '0';
                        hold_seg_2     <=  '1';
                        hold_seg_3     <=  '1';
                        hold_seg_4     <=  '1';
                        hold_seg_5     <=  '1';
                        hold_seg_6     <=  '1';
                        hold_seg_7     <=  '1';
                        in_ctrl_all_cb <=  '1';
                        hold_all_out   <=  '0';
                        in_ctrl_all_out<=  '0';
                        counter_en     <=  '0';
                        currentstate   <= state_3;					
                    WHEN state_3		 =>
                        hold_all_in    <=  '1';
                        hold_buf_3     <=  '1';
                        hold_buf_2     <=  '1';
                        hold_buf_1     <=  '0';
                        in_ctrl_buf_3  <=  '0';
                        in_ctrl_buf_2  <=  '0';
                        in_ctrl_buf_1  <=  '1';
                        pos_hold_ctrl  <=  '1';
                        Shuf_Ctrl_1    <=  "000";
                        Shuf_Ctrl_2    <=  "001";
                        Shuf_Ctrl_3    <=  "000";
                        Shuf_Ctrl_4    <=  "010";
                        Shuf_Ctrl_5    <=  "000";
                        Shuf_Ctrl_6    <=  "011";
                        Shuf_Ctrl_7    <=  "000";
                        Shuf_Ctrl_8    <=  "100";
                        Type_Sel_1     <=  "000";
                        Type_Sel_2     <=  "001";
                        Type_Sel_3     <=  "000";
                        Type_Sel_4     <=  "001";
                        Type_Sel_5     <=  "000";
                        Type_Sel_6     <=  "001";
                        Type_Sel_7     <=  "000";
                        Type_Sel_8     <=  "001";
                        Bypass_Sel_0   <=  "000";
                        Bypass_Sel_1   <=  "000";
                        Bypass_Sel_2   <=  "000";
                        Bypass_Sel_3   <=  "000";
                        Bypass_Sel_4   <=  "000";
                        Bypass_Sel_5   <=  "000";
                        Bypass_Sel_6   <=  "000";
                        Bypass_Sel_7   <=  "000";
                        DeShuf_Ctrl_0  <=  "000";
                        DeShuf_Ctrl_1  <=  "001";
                        DeShuf_Ctrl_2  <=  "011";
                        DeShuf_Ctrl_3  <=  "101";
                        DeShuf_Ctrl_4  <=  "111";
                        DeShuf_Ctrl_5  <=  "000";
                        DeShuf_Ctrl_6  <=  "000";
                        DeShuf_Ctrl_7  <=  "000";
                        Bypass_EN_0    <=  '1';
                        Bypass_EN_1    <=  '0';
                        Bypass_EN_2    <=  '0';
                        Bypass_EN_3    <=  '0';
                        Bypass_EN_4    <=  '0';
                        Bypass_EN_5    <=  '0';
                        Bypass_EN_6    <=  '0';
                        Bypass_EN_7    <=  '0';
                        Hold_Ctrl_0    <=  '0';
                        Hold_Ctrl_1    <=  '0';
                        Hold_Ctrl_2    <=  '0';
                        Hold_Ctrl_3    <=  '0';
                        Hold_Ctrl_4    <=  '0';
                        Hold_Ctrl_5    <=  '0';
                        Hold_Ctrl_6    <=  '0';
                        Hold_Ctrl_7    <=  '0';
                        DFF_Ctrl_0     <=  '0';
                        DFF_Ctrl_1     <=  '0';
                        DFF_Ctrl_2     <=  '0';
                        DFF_Ctrl_3     <=  '0';
                        DFF_Ctrl_4     <=  '0';
                        DFF_Ctrl_5     <=  '0';
                        DFF_Ctrl_6     <=  '0';
                        DFF_Ctrl_7     <=  '0';
                        hold_seg_0     <=  '1';
                        hold_seg_1     <=  '1';
                        hold_seg_2     <=  '1';
                        hold_seg_3     <=  '1';
                        hold_seg_4     <=  '1';
                        hold_seg_5     <=  '1';
                        hold_seg_6     <=  '1';
                        hold_seg_7     <=  '1';
                        in_ctrl_all_cb <=  '1';
                        hold_all_out   <=  '0';
                        in_ctrl_all_out<=  '0';
                        counter_en     <=  '0';
                        currentstate   <= state_4;					
                    WHEN state_4		 =>
                        hold_all_in    <=  '0';
                        hold_buf_3     <=  '1';
                        hold_buf_2     <=  '1';
                        hold_buf_1     <=  '0';
                        in_ctrl_buf_3  <=  '0';
                        in_ctrl_buf_2  <=  '0';
                        in_ctrl_buf_1  <=  '1';
                        pos_hold_ctrl  <=  '1';
                        Shuf_Ctrl_1    <=  "000";
                        Shuf_Ctrl_2    <=  "111";
                        Shuf_Ctrl_3    <=  "000";
                        Shuf_Ctrl_4    <=  "110";
                        Shuf_Ctrl_5    <=  "000";
                        Shuf_Ctrl_6    <=  "101";
                        Shuf_Ctrl_7    <=  "000";
                        Shuf_Ctrl_8    <=  "000";
                        Type_Sel_1     <=  "000";
                        Type_Sel_2     <=  "101";
                        Type_Sel_3     <=  "000";
                        Type_Sel_4     <=  "101";
                        Type_Sel_5     <=  "000";
                        Type_Sel_6     <=  "101";
                        Type_Sel_7     <=  "000";
                        Type_Sel_8     <=  "000";
                        Bypass_Sel_0   <=  "000";
                        Bypass_Sel_1   <=  "000";
                        Bypass_Sel_2   <=  "000";
                        Bypass_Sel_3   <=  "000";
                        Bypass_Sel_4   <=  "000";
                        Bypass_Sel_5   <=  "000";
                        Bypass_Sel_6   <=  "000";
                        Bypass_Sel_7   <=  "000";
                        DeShuf_Ctrl_0  <=  "000";
                        DeShuf_Ctrl_1  <=  "000";
                        DeShuf_Ctrl_2  <=  "000";
                        DeShuf_Ctrl_3  <=  "000";
                        DeShuf_Ctrl_4  <=  "000";
                        DeShuf_Ctrl_5  <=  "101";
                        DeShuf_Ctrl_6  <=  "011";
                        DeShuf_Ctrl_7  <=  "001";
                        Bypass_EN_0    <=  '1';
                        Bypass_EN_1    <=  '0';
                        Bypass_EN_2    <=  '0';
                        Bypass_EN_3    <=  '0';
                        Bypass_EN_4    <=  '0';
                        Bypass_EN_5    <=  '0';
                        Bypass_EN_6    <=  '0';
                        Bypass_EN_7    <=  '0';
                        Hold_Ctrl_0    <=  '1';
                        Hold_Ctrl_1    <=  '1';
                        Hold_Ctrl_2    <=  '1';
                        Hold_Ctrl_3    <=  '1';
                        Hold_Ctrl_4    <=  '1';
                        Hold_Ctrl_5    <=  '0';
                        Hold_Ctrl_6    <=  '0';
                        Hold_Ctrl_7    <=  '0';
                        DFF_Ctrl_0     <=  '1';
                        DFF_Ctrl_1     <=  '1';
                        DFF_Ctrl_2     <=  '1';
                        DFF_Ctrl_3     <=  '1';
                        DFF_Ctrl_4     <=  '1';
                        DFF_Ctrl_5     <=  '0';
                        DFF_Ctrl_6     <=  '0';
                        DFF_Ctrl_7     <=  '0';
                        hold_seg_0     <=  '1';
                        hold_seg_1     <=  '1';
                        hold_seg_2     <=  '0';
                        hold_seg_3     <=  '1';
                        hold_seg_4     <=  '1';
                        hold_seg_5     <=  '1';
                        hold_seg_6     <=  '1';
                        hold_seg_7     <=  '1';
                        in_ctrl_all_cb <=  '1';
                        hold_all_out   <=  '0';
                        in_ctrl_all_out<=  '0';
                        counter_en     <=  '0';
                        currentstate   <= state_5;					
                    WHEN state_5		 =>
                        hold_all_in    <=  '0';
                        hold_buf_3     <=  '1';
                        hold_buf_2     <=  '1';
                        hold_buf_1     <=  '0';
                        in_ctrl_buf_3  <=  '0';
                        in_ctrl_buf_2  <=  '0';
                        in_ctrl_buf_1  <=  '1';
                        pos_hold_ctrl  <=  '1';
                        Shuf_Ctrl_1    <=  "101";
                        Shuf_Ctrl_2    <=  "110";
                        Shuf_Ctrl_3    <=  "001";
                        Shuf_Ctrl_4    <=  "100";
                        Shuf_Ctrl_5    <=  "111";
                        Shuf_Ctrl_6    <=  "010";
                        Shuf_Ctrl_7    <=  "011";
                        Shuf_Ctrl_8    <=  "000";
                        Type_Sel_1     <=  "101";
                        Type_Sel_2     <=  "111";
                        Type_Sel_3     <=  "001";
                        Type_Sel_4     <=  "101";
                        Type_Sel_5     <=  "111";
                        Type_Sel_6     <=  "001";
                        Type_Sel_7     <=  "101";
                        Type_Sel_8     <=  "000";
                        Bypass_Sel_0   <=  "000";
                        Bypass_Sel_1   <=  "000";
                        Bypass_Sel_2   <=  "000";
                        Bypass_Sel_3   <=  "000";
                        Bypass_Sel_4   <=  "000";
                        Bypass_Sel_5   <=  "000";
                        Bypass_Sel_6   <=  "000";
                        Bypass_Sel_7   <=  "000";
                        DeShuf_Ctrl_0  <=  "000";
                        DeShuf_Ctrl_1  <=  "010";
                        DeShuf_Ctrl_2  <=  "101";
                        DeShuf_Ctrl_3  <=  "110";
                        DeShuf_Ctrl_4  <=  "011";
                        DeShuf_Ctrl_5  <=  "000";
                        DeShuf_Ctrl_6  <=  "001";
                        DeShuf_Ctrl_7  <=  "100";
                        Bypass_EN_0    <=  '1';
                        Bypass_EN_1    <=  '0';
                        Bypass_EN_2    <=  '0';
                        Bypass_EN_3    <=  '0';
                        Bypass_EN_4    <=  '0';
                        Bypass_EN_5    <=  '0';
                        Bypass_EN_6    <=  '0';
                        Bypass_EN_7    <=  '0';
                        Hold_Ctrl_0    <=  '0';
                        Hold_Ctrl_1    <=  '0';
                        Hold_Ctrl_2    <=  '0';
                        Hold_Ctrl_3    <=  '0';
                        Hold_Ctrl_4    <=  '0';
                        Hold_Ctrl_5    <=  '0';
                        Hold_Ctrl_6    <=  '0';
                        Hold_Ctrl_7    <=  '0';
                        DFF_Ctrl_0     <=  '0';
                        DFF_Ctrl_1     <=  '0';
                        DFF_Ctrl_2     <=  '0';
                        DFF_Ctrl_3     <=  '0';
                        DFF_Ctrl_4     <=  '0';
                        DFF_Ctrl_5     <=  '0';
                        DFF_Ctrl_6     <=  '0';
                        DFF_Ctrl_7     <=  '0';
                        hold_seg_0     <=  '1';
                        hold_seg_1     <=  '1';
                        hold_seg_2     <=  '1';
                        hold_seg_3     <=  '0';
                        hold_seg_4     <=  '1';
                        hold_seg_5     <=  '1';
                        hold_seg_6     <=  '1';
                        hold_seg_7     <=  '1';
                        in_ctrl_all_cb <=  '1';
                        hold_all_out   <=  '0';
                        in_ctrl_all_out<=  '0';
                        counter_en     <=  '0';
                        currentstate   <= state_6;					
                    WHEN state_6		 =>
                        hold_all_in    <=  '1';
                        hold_buf_3     <=  '1';
                        hold_buf_2     <=  '0';
                        hold_buf_1     <=  '1';
                        in_ctrl_buf_3  <=  '0';
                        in_ctrl_buf_2  <=  '1';
                        in_ctrl_buf_1  <=  '0';
                        pos_hold_ctrl  <=  '1';
                        Shuf_Ctrl_1    <=  "000";
                        Shuf_Ctrl_2    <=  "000";
                        Shuf_Ctrl_3    <=  "000";
                        Shuf_Ctrl_4    <=  "001";
                        Shuf_Ctrl_5    <=  "000";
                        Shuf_Ctrl_6    <=  "000";
                        Shuf_Ctrl_7    <=  "000";
                        Shuf_Ctrl_8    <=  "010";
                        Type_Sel_1     <=  "000";
                        Type_Sel_2     <=  "000";
                        Type_Sel_3     <=  "000";
                        Type_Sel_4     <=  "001";
                        Type_Sel_5     <=  "000";
                        Type_Sel_6     <=  "000";
                        Type_Sel_7     <=  "000";
                        Type_Sel_8     <=  "001";
                        Bypass_Sel_0   <=  "000";
                        Bypass_Sel_1   <=  "000";
                        Bypass_Sel_2   <=  "000";
                        Bypass_Sel_3   <=  "000";
                        Bypass_Sel_4   <=  "101";
                        Bypass_Sel_5   <=  "000";
                        Bypass_Sel_6   <=  "000";
                        Bypass_Sel_7   <=  "000";
                        DeShuf_Ctrl_0  <=  "000";
                        DeShuf_Ctrl_1  <=  "011";
                        DeShuf_Ctrl_2  <=  "111";
                        DeShuf_Ctrl_3  <=  "000";
                        DeShuf_Ctrl_4  <=  "000";
                        DeShuf_Ctrl_5  <=  "000";
                        DeShuf_Ctrl_6  <=  "000";
                        DeShuf_Ctrl_7  <=  "000";
                        Bypass_EN_0    <=  '1';
                        Bypass_EN_1    <=  '0';
                        Bypass_EN_2    <=  '0';
                        Bypass_EN_3    <=  '0';
                        Bypass_EN_4    <=  '1';
                        Bypass_EN_5    <=  '0';
                        Bypass_EN_6    <=  '0';
                        Bypass_EN_7    <=  '0';
                        Hold_Ctrl_0    <=  '0';
                        Hold_Ctrl_1    <=  '0';
                        Hold_Ctrl_2    <=  '0';
                        Hold_Ctrl_3    <=  '0';
                        Hold_Ctrl_4    <=  '0';
                        Hold_Ctrl_5    <=  '0';
                        Hold_Ctrl_6    <=  '0';
                        Hold_Ctrl_7    <=  '0';
                        DFF_Ctrl_0     <=  '0';
                        DFF_Ctrl_1     <=  '0';
                        DFF_Ctrl_2     <=  '0';
                        DFF_Ctrl_3     <=  '0';
                        DFF_Ctrl_4     <=  '0';
                        DFF_Ctrl_5     <=  '0';
                        DFF_Ctrl_6     <=  '0';
                        DFF_Ctrl_7     <=  '0';
                        hold_seg_0     <=  '1';
                        hold_seg_1     <=  '1';
                        hold_seg_2     <=  '1';
                        hold_seg_3     <=  '1';
                        hold_seg_4     <=  '1';
                        hold_seg_5     <=  '1';
                        hold_seg_6     <=  '1';
                        hold_seg_7     <=  '1';
                        in_ctrl_all_cb <=  '1';
                        hold_all_out   <=  '0';
                        in_ctrl_all_out<=  '0';
                        counter_en     <=  '0';
                        currentstate   <= state_7;					
                    WHEN state_7		 =>
                        hold_all_in    <=  '1';
                        hold_buf_3     <=  '0';
                        hold_buf_2     <=  '1';
                        hold_buf_1     <=  '1';
                        in_ctrl_buf_3  <=  '1';
                        in_ctrl_buf_2  <=  '0';
                        in_ctrl_buf_1  <=  '0';
                        pos_hold_ctrl  <=  '1';
                        Shuf_Ctrl_1    <=  "000";
                        Shuf_Ctrl_2    <=  "000";
                        Shuf_Ctrl_3    <=  "000";
                        Shuf_Ctrl_4    <=  "011";
                        Shuf_Ctrl_5    <=  "000";
                        Shuf_Ctrl_6    <=  "000";
                        Shuf_Ctrl_7    <=  "000";
                        Shuf_Ctrl_8    <=  "000";
                        Type_Sel_1     <=  "000";
                        Type_Sel_2     <=  "000";
                        Type_Sel_3     <=  "000";
                        Type_Sel_4     <=  "101";
                        Type_Sel_5     <=  "000";
                        Type_Sel_6     <=  "000";
                        Type_Sel_7     <=  "000";
                        Type_Sel_8     <=  "000";
                        Bypass_Sel_0   <=  "000";
                        Bypass_Sel_1   <=  "000";
                        Bypass_Sel_2   <=  "000";
                        Bypass_Sel_3   <=  "000";
                        Bypass_Sel_4   <=  "000";
                        Bypass_Sel_5   <=  "000";
                        Bypass_Sel_6   <=  "000";
                        Bypass_Sel_7   <=  "000";
                        DeShuf_Ctrl_0  <=  "000";
                        DeShuf_Ctrl_1  <=  "000";
                        DeShuf_Ctrl_2  <=  "000";
                        DeShuf_Ctrl_3  <=  "011";
                        DeShuf_Ctrl_4  <=  "000";
                        DeShuf_Ctrl_5  <=  "000";
                        DeShuf_Ctrl_6  <=  "000";
                        DeShuf_Ctrl_7  <=  "000";
                        Bypass_EN_0    <=  '1';
                        Bypass_EN_1    <=  '0';
                        Bypass_EN_2    <=  '0';
                        Bypass_EN_3    <=  '0';
                        Bypass_EN_4    <=  '0';
                        Bypass_EN_5    <=  '0';
                        Bypass_EN_6    <=  '0';
                        Bypass_EN_7    <=  '0';
                        Hold_Ctrl_0    <=  '1';
                        Hold_Ctrl_1    <=  '1';
                        Hold_Ctrl_2    <=  '1';
                        Hold_Ctrl_3    <=  '0';
                        Hold_Ctrl_4    <=  '1';
                        Hold_Ctrl_5    <=  '0';
                        Hold_Ctrl_6    <=  '0';
                        Hold_Ctrl_7    <=  '0';
                        DFF_Ctrl_0     <=  '1';
                        DFF_Ctrl_1     <=  '1';
                        DFF_Ctrl_2     <=  '1';
                        DFF_Ctrl_3     <=  '0';
                        DFF_Ctrl_4     <=  '1';
                        DFF_Ctrl_5     <=  '0';
                        DFF_Ctrl_6     <=  '0';
                        DFF_Ctrl_7     <=  '0';
                        hold_seg_0     <=  '1';
                        hold_seg_1     <=  '1';
                        hold_seg_2     <=  '1';
                        hold_seg_3     <=  '1';
                        hold_seg_4     <=  '1';
                        hold_seg_5     <=  '1';
                        hold_seg_6     <=  '1';
                        hold_seg_7     <=  '1';
                        in_ctrl_all_cb <=  '1';
                        hold_all_out   <=  '0';
                        in_ctrl_all_out<=  '0';
                        counter_en     <=  '0';
                        currentstate   <= state_8;					
                    WHEN state_8		 =>
                        hold_all_in    <=  '1';
                        hold_buf_3     <=  '1';
                        hold_buf_2     <=  '1';
                        hold_buf_1     <=  '1';
                        in_ctrl_buf_3  <=  '0';
                        in_ctrl_buf_2  <=  '0';
                        in_ctrl_buf_1  <=  '0';
                        pos_hold_ctrl  <=  '1';
                        Shuf_Ctrl_1    <=  "000";
                        Shuf_Ctrl_2    <=  "000";
                        Shuf_Ctrl_3    <=  "000";
                        Shuf_Ctrl_4    <=  "101";
                        Shuf_Ctrl_5    <=  "000";
                        Shuf_Ctrl_6    <=  "000";
                        Shuf_Ctrl_7    <=  "000";
                        Shuf_Ctrl_8    <=  "110";
                        Type_Sel_1     <=  "000";
                        Type_Sel_2     <=  "000";
                        Type_Sel_3     <=  "000";
                        Type_Sel_4     <=  "111";
                        Type_Sel_5     <=  "000";
                        Type_Sel_6     <=  "000";
                        Type_Sel_7     <=  "000";
                        Type_Sel_8     <=  "111";
                        Bypass_Sel_0   <=  "000";
                        Bypass_Sel_1   <=  "000";
                        Bypass_Sel_2   <=  "000";
                        Bypass_Sel_3   <=  "000";
                        Bypass_Sel_4   <=  "000";
                        Bypass_Sel_5   <=  "000";
                        Bypass_Sel_6   <=  "000";
                        Bypass_Sel_7   <=  "000";
                        DeShuf_Ctrl_0  <=  "000";
                        DeShuf_Ctrl_1  <=  "000";
                        DeShuf_Ctrl_2  <=  "000";
                        DeShuf_Ctrl_3  <=  "000";
                        DeShuf_Ctrl_4  <=  "000";
                        DeShuf_Ctrl_5  <=  "011";
                        DeShuf_Ctrl_6  <=  "111";
                        DeShuf_Ctrl_7  <=  "000";
                        Bypass_EN_0    <=  '1';
                        Bypass_EN_1    <=  '0';
                        Bypass_EN_2    <=  '0';
                        Bypass_EN_3    <=  '0';
                        Bypass_EN_4    <=  '0';
                        Bypass_EN_5    <=  '0';
                        Bypass_EN_6    <=  '0';
                        Bypass_EN_7    <=  '0';
                        Hold_Ctrl_0    <=  '1';
                        Hold_Ctrl_1    <=  '1';
                        Hold_Ctrl_2    <=  '1';
                        Hold_Ctrl_3    <=  '1';
                        Hold_Ctrl_4    <=  '1';
                        Hold_Ctrl_5    <=  '0';
                        Hold_Ctrl_6    <=  '0';
                        Hold_Ctrl_7    <=  '0';
                        DFF_Ctrl_0     <=  '1';
                        DFF_Ctrl_1     <=  '1';
                        DFF_Ctrl_2     <=  '1';
                        DFF_Ctrl_3     <=  '1';
                        DFF_Ctrl_4     <=  '1';
                        DFF_Ctrl_5     <=  '0';
                        DFF_Ctrl_6     <=  '0';
                        DFF_Ctrl_7     <=  '0';
                        hold_seg_0     <=  '1';
                        hold_seg_1     <=  '1';
                        hold_seg_2     <=  '1';
                        hold_seg_3     <=  '1';
                        hold_seg_4     <=  '1';
                        hold_seg_5     <=  '1';
                        hold_seg_6     <=  '1';
                        hold_seg_7     <=  '1';
                        in_ctrl_all_cb <=  '1';
                        hold_all_out   <=  '0';
                        in_ctrl_all_out<=  '0';
                        counter_en     <=  '0';
                        currentstate   <= state_9;					
                    WHEN state_9		 =>
                        hold_all_in    <=  '0';
                        hold_buf_3     <=  '0';
                        hold_buf_2     <=  '0';
                        hold_buf_1     <=  '0';
                        in_ctrl_buf_3  <=  '0';
                        in_ctrl_buf_2  <=  '0';
                        in_ctrl_buf_1  <=  '0';
                        pos_hold_ctrl  <=  '1';
                        Shuf_Ctrl_1    <=  "000";
                        Shuf_Ctrl_2    <=  "000";
                        Shuf_Ctrl_3    <=  "000";
                        Shuf_Ctrl_4    <=  "111";
                        Shuf_Ctrl_5    <=  "000";
                        Shuf_Ctrl_6    <=  "000";
                        Shuf_Ctrl_7    <=  "000";
                        Shuf_Ctrl_8    <=  "000";
                        Type_Sel_1     <=  "000";
                        Type_Sel_2     <=  "000";
                        Type_Sel_3     <=  "000";
                        Type_Sel_4     <=  "011";
                        Type_Sel_5     <=  "000";
                        Type_Sel_6     <=  "000";
                        Type_Sel_7     <=  "000";
                        Type_Sel_8     <=  "000";
                        Bypass_Sel_0   <=  "000";
                        Bypass_Sel_1   <=  "000";
                        Bypass_Sel_2   <=  "000";
                        Bypass_Sel_3   <=  "000";
                        Bypass_Sel_4   <=  "000";
                        Bypass_Sel_5   <=  "000";
                        Bypass_Sel_6   <=  "000";
                        Bypass_Sel_7   <=  "000";
                        DeShuf_Ctrl_0  <=  "000";
                        DeShuf_Ctrl_1  <=  "000";
                        DeShuf_Ctrl_2  <=  "000";
                        DeShuf_Ctrl_3  <=  "000";
                        DeShuf_Ctrl_4  <=  "000";
                        DeShuf_Ctrl_5  <=  "000";
                        DeShuf_Ctrl_6  <=  "000";
                        DeShuf_Ctrl_7  <=  "011";
                        Bypass_EN_0    <=  '1';
                        Bypass_EN_1    <=  '0';
                        Bypass_EN_2    <=  '0';
                        Bypass_EN_3    <=  '0';
                        Bypass_EN_4    <=  '0';
                        Bypass_EN_5    <=  '0';
                        Bypass_EN_6    <=  '0';
                        Bypass_EN_7    <=  '0';
                        Hold_Ctrl_0    <=  '1';
                        Hold_Ctrl_1    <=  '1';
                        Hold_Ctrl_2    <=  '1';
                        Hold_Ctrl_3    <=  '1';
                        Hold_Ctrl_4    <=  '1';
                        Hold_Ctrl_5    <=  '1';
                        Hold_Ctrl_6    <=  '1';
                        Hold_Ctrl_7    <=  '0';
                        DFF_Ctrl_0     <=  '1';
                        DFF_Ctrl_1     <=  '1';
                        DFF_Ctrl_2     <=  '1';
                        DFF_Ctrl_3     <=  '1';
                        DFF_Ctrl_4     <=  '1';
                        DFF_Ctrl_5     <=  '1';
                        DFF_Ctrl_6     <=  '1';
                        DFF_Ctrl_7     <=  '0';
                        hold_seg_0     <=  '1';
                        hold_seg_1     <=  '1';
                        hold_seg_2     <=  '1';
                        hold_seg_3     <=  '1';
                        hold_seg_4     <=  '0';
                        hold_seg_5     <=  '1';
                        hold_seg_6     <=  '1';
                        hold_seg_7     <=  '1';
                        in_ctrl_all_cb <=  '1';
                        hold_all_out   <=  '0';
                        in_ctrl_all_out<=  '0';
                        counter_en     <=  '0';
                        currentstate   <= state_10;					
                    WHEN state_10		 =>
                        hold_all_in    <=  '0';
                        hold_buf_3     <=  '0';
                        hold_buf_2     <=  '0';
                        hold_buf_1     <=  '0';
                        in_ctrl_buf_3  <=  '0';
                        in_ctrl_buf_2  <=  '0';
                        in_ctrl_buf_1  <=  '0';
                        pos_hold_ctrl  <=  '1';
                        Shuf_Ctrl_1    <=  "011";
                        Shuf_Ctrl_2    <=  "110";
                        Shuf_Ctrl_3    <=  "111";
                        Shuf_Ctrl_4    <=  "100";
                        Shuf_Ctrl_5    <=  "001";
                        Shuf_Ctrl_6    <=  "010";
                        Shuf_Ctrl_7    <=  "101";
                        Shuf_Ctrl_8    <=  "000";
                        Type_Sel_1     <=  "101";
                        Type_Sel_2     <=  "011";
                        Type_Sel_3     <=  "010";
                        Type_Sel_4     <=  "111";
                        Type_Sel_5     <=  "001";
                        Type_Sel_6     <=  "101";
                        Type_Sel_7     <=  "011";
                        Type_Sel_8     <=  "000";
                        Bypass_Sel_0   <=  "000";
                        Bypass_Sel_1   <=  "000";
                        Bypass_Sel_2   <=  "000";
                        Bypass_Sel_3   <=  "000";
                        Bypass_Sel_4   <=  "000";
                        Bypass_Sel_5   <=  "000";
                        Bypass_Sel_6   <=  "000";
                        Bypass_Sel_7   <=  "000";
                        DeShuf_Ctrl_0  <=  "000";
                        DeShuf_Ctrl_1  <=  "100";
                        DeShuf_Ctrl_2  <=  "101";
                        DeShuf_Ctrl_3  <=  "000";
                        DeShuf_Ctrl_4  <=  "011";
                        DeShuf_Ctrl_5  <=  "110";
                        DeShuf_Ctrl_6  <=  "001";
                        DeShuf_Ctrl_7  <=  "010";
                        Bypass_EN_0    <=  '1';
                        Bypass_EN_1    <=  '0';
                        Bypass_EN_2    <=  '0';
                        Bypass_EN_3    <=  '0';
                        Bypass_EN_4    <=  '0';
                        Bypass_EN_5    <=  '0';
                        Bypass_EN_6    <=  '0';
                        Bypass_EN_7    <=  '0';
                        Hold_Ctrl_0    <=  '0';
                        Hold_Ctrl_1    <=  '0';
                        Hold_Ctrl_2    <=  '0';
                        Hold_Ctrl_3    <=  '0';
                        Hold_Ctrl_4    <=  '0';
                        Hold_Ctrl_5    <=  '0';
                        Hold_Ctrl_6    <=  '0';
                        Hold_Ctrl_7    <=  '0';
                        DFF_Ctrl_0     <=  '0';
                        DFF_Ctrl_1     <=  '0';
                        DFF_Ctrl_2     <=  '0';
                        DFF_Ctrl_3     <=  '0';
                        DFF_Ctrl_4     <=  '0';
                        DFF_Ctrl_5     <=  '0';
                        DFF_Ctrl_6     <=  '0';
                        DFF_Ctrl_7     <=  '0';
                        hold_seg_0     <=  '1';
                        hold_seg_1     <=  '1';
                        hold_seg_2     <=  '1';
                        hold_seg_3     <=  '1';
                        hold_seg_4     <=  '1';
                        hold_seg_5     <=  '0';
                        hold_seg_6     <=  '1';
                        hold_seg_7     <=  '1';
                        in_ctrl_all_cb <=  '1';
                        hold_all_out   <=  '0';
                        in_ctrl_all_out<=  '0';
                        counter_en     <=  '0';
                        currentstate   <= state_11;					
                    WHEN state_11		 =>
                        hold_all_in    <=  '1';
                        hold_buf_3     <=  '1';
                        hold_buf_2     <=  '1';
                        hold_buf_1     <=  '1';
                        in_ctrl_buf_3  <=  '0';
                        in_ctrl_buf_2  <=  '0';
                        in_ctrl_buf_1  <=  '0';
                        pos_hold_ctrl  <=  '1';
                        Shuf_Ctrl_1    <=  "000";
                        Shuf_Ctrl_2    <=  "011";
                        Shuf_Ctrl_3    <=  "000";
                        Shuf_Ctrl_4    <=  "010";
                        Shuf_Ctrl_5    <=  "000";
                        Shuf_Ctrl_6    <=  "001";
                        Shuf_Ctrl_7    <=  "000";
                        Shuf_Ctrl_8    <=  "100";
                        Type_Sel_1     <=  "000";
                        Type_Sel_2     <=  "111";
                        Type_Sel_3     <=  "000";
                        Type_Sel_4     <=  "101";
                        Type_Sel_5     <=  "000";
                        Type_Sel_6     <=  "001";
                        Type_Sel_7     <=  "000";
                        Type_Sel_8     <=  "111";
                        Bypass_Sel_0   <=  "000";
                        Bypass_Sel_1   <=  "000";
                        Bypass_Sel_2   <=  "000";
                        Bypass_Sel_3   <=  "000";
                        Bypass_Sel_4   <=  "000";
                        Bypass_Sel_5   <=  "000";
                        Bypass_Sel_6   <=  "000";
                        Bypass_Sel_7   <=  "000";
                        DeShuf_Ctrl_0  <=  "000";
                        DeShuf_Ctrl_1  <=  "101";
                        DeShuf_Ctrl_2  <=  "011";
                        DeShuf_Ctrl_3  <=  "001";
                        DeShuf_Ctrl_4  <=  "111";
                        DeShuf_Ctrl_5  <=  "000";
                        DeShuf_Ctrl_6  <=  "000";
                        DeShuf_Ctrl_7  <=  "000";
                        Bypass_EN_0    <=  '1';
                        Bypass_EN_1    <=  '0';
                        Bypass_EN_2    <=  '0';
                        Bypass_EN_3    <=  '0';
                        Bypass_EN_4    <=  '0';
                        Bypass_EN_5    <=  '0';
                        Bypass_EN_6    <=  '0';
                        Bypass_EN_7    <=  '0';
                        Hold_Ctrl_0    <=  '0';
                        Hold_Ctrl_1    <=  '0';
                        Hold_Ctrl_2    <=  '0';
                        Hold_Ctrl_3    <=  '0';
                        Hold_Ctrl_4    <=  '0';
                        Hold_Ctrl_5    <=  '0';
                        Hold_Ctrl_6    <=  '0';
                        Hold_Ctrl_7    <=  '0';
                        DFF_Ctrl_0     <=  '0';
                        DFF_Ctrl_1     <=  '0';
                        DFF_Ctrl_2     <=  '0';
                        DFF_Ctrl_3     <=  '0';
                        DFF_Ctrl_4     <=  '0';
                        DFF_Ctrl_5     <=  '0';
                        DFF_Ctrl_6     <=  '0';
                        DFF_Ctrl_7     <=  '0';
                        hold_seg_0     <=  '1';
                        hold_seg_1     <=  '1';
                        hold_seg_2     <=  '1';
                        hold_seg_3     <=  '1';
                        hold_seg_4     <=  '1';
                        hold_seg_5     <=  '1';
                        hold_seg_6     <=  '1';
                        hold_seg_7     <=  '1';
                        in_ctrl_all_cb <=  '1';
                        hold_all_out   <=  '0';
                        in_ctrl_all_out<=  '0';
                        counter_en     <=  '0';
                        currentstate   <= state_12;					
                    WHEN state_12		 =>
                        hold_all_in    <=  '0';
                        hold_buf_3     <=  '0';
                        hold_buf_2     <=  '0';
                        hold_buf_1     <=  '0';
                        in_ctrl_buf_3  <=  '0';
                        in_ctrl_buf_2  <=  '0';
                        in_ctrl_buf_1  <=  '0';
                        pos_hold_ctrl  <=  '1';
                        Shuf_Ctrl_1    <=  "000";
                        Shuf_Ctrl_2    <=  "101";
                        Shuf_Ctrl_3    <=  "000";
                        Shuf_Ctrl_4    <=  "110";
                        Shuf_Ctrl_5    <=  "000";
                        Shuf_Ctrl_6    <=  "111";
                        Shuf_Ctrl_7    <=  "000";
                        Shuf_Ctrl_8    <=  "000";
                        Type_Sel_1     <=  "000";
                        Type_Sel_2     <=  "011";
                        Type_Sel_3     <=  "000";
                        Type_Sel_4     <=  "010";
                        Type_Sel_5     <=  "000";
                        Type_Sel_6     <=  "110";
                        Type_Sel_7     <=  "000";
                        Type_Sel_8     <=  "000";
                        Bypass_Sel_0   <=  "000";
                        Bypass_Sel_1   <=  "000";
                        Bypass_Sel_2   <=  "000";
                        Bypass_Sel_3   <=  "000";
                        Bypass_Sel_4   <=  "000";
                        Bypass_Sel_5   <=  "000";
                        Bypass_Sel_6   <=  "000";
                        Bypass_Sel_7   <=  "000";
                        DeShuf_Ctrl_0  <=  "000";
                        DeShuf_Ctrl_1  <=  "000";
                        DeShuf_Ctrl_2  <=  "000";
                        DeShuf_Ctrl_3  <=  "000";
                        DeShuf_Ctrl_4  <=  "000";
                        DeShuf_Ctrl_5  <=  "001";
                        DeShuf_Ctrl_6  <=  "011";
                        DeShuf_Ctrl_7  <=  "101";
                        Bypass_EN_0    <=  '1';
                        Bypass_EN_1    <=  '0';
                        Bypass_EN_2    <=  '0';
                        Bypass_EN_3    <=  '0';
                        Bypass_EN_4    <=  '0';
                        Bypass_EN_5    <=  '0';
                        Bypass_EN_6    <=  '0';
                        Bypass_EN_7    <=  '0';
                        Hold_Ctrl_0    <=  '1';
                        Hold_Ctrl_1    <=  '1';
                        Hold_Ctrl_2    <=  '1';
                        Hold_Ctrl_3    <=  '1';
                        Hold_Ctrl_4    <=  '1';
                        Hold_Ctrl_5    <=  '0';
                        Hold_Ctrl_6    <=  '0';
                        Hold_Ctrl_7    <=  '0';
                        DFF_Ctrl_0     <=  '1';
                        DFF_Ctrl_1     <=  '1';
                        DFF_Ctrl_2     <=  '1';
                        DFF_Ctrl_3     <=  '1';
                        DFF_Ctrl_4     <=  '1';
                        DFF_Ctrl_5     <=  '0';
                        DFF_Ctrl_6     <=  '0';
                        DFF_Ctrl_7     <=  '0';
                        hold_seg_0     <=  '1';
                        hold_seg_1     <=  '1';
                        hold_seg_2     <=  '1';
                        hold_seg_3     <=  '1';
                        hold_seg_4     <=  '1';
                        hold_seg_5     <=  '1';
                        hold_seg_6     <=  '0';
                        hold_seg_7     <=  '1';
                        in_ctrl_all_cb <=  '1';
                        hold_all_out   <=  '0';
                        in_ctrl_all_out<=  '0';
                        counter_en     <=  '0';
                        currentstate   <= state_13;					
                    WHEN state_13		 =>
                        hold_all_in    <=  '0';
                        hold_buf_3     <=  '1';
                        hold_buf_2     <=  '1';
                        hold_buf_1     <=  '1';
                        in_ctrl_buf_3  <=  '0';
                        in_ctrl_buf_2  <=  '0';
                        in_ctrl_buf_1  <=  '0';
                        pos_hold_ctrl  <=  '0';
                        Shuf_Ctrl_1    <=  "111";
                        Shuf_Ctrl_2    <=  "010";
                        Shuf_Ctrl_3    <=  "101";
                        Shuf_Ctrl_4    <=  "100";
                        Shuf_Ctrl_5    <=  "011";
                        Shuf_Ctrl_6    <=  "110";
                        Shuf_Ctrl_7    <=  "001";
                        Shuf_Ctrl_8    <=  "000";
                        Type_Sel_1     <=  "100";
                        Type_Sel_2     <=  "101";
                        Type_Sel_3     <=  "010";
                        Type_Sel_4     <=  "011";
                        Type_Sel_5     <=  "111";
                        Type_Sel_6     <=  "110";
                        Type_Sel_7     <=  "001";
                        Type_Sel_8     <=  "000";
                        Bypass_Sel_0   <=  "000";
                        Bypass_Sel_1   <=  "000";
                        Bypass_Sel_2   <=  "000";
                        Bypass_Sel_3   <=  "000";
                        Bypass_Sel_4   <=  "000";
                        Bypass_Sel_5   <=  "000";
                        Bypass_Sel_6   <=  "000";
                        Bypass_Sel_7   <=  "000";
                        DeShuf_Ctrl_0  <=  "000";
                        DeShuf_Ctrl_1  <=  "110";
                        DeShuf_Ctrl_2  <=  "001";
                        DeShuf_Ctrl_3  <=  "100";
                        DeShuf_Ctrl_4  <=  "011";
                        DeShuf_Ctrl_5  <=  "010";
                        DeShuf_Ctrl_6  <=  "101";
                        DeShuf_Ctrl_7  <=  "000";
                        Bypass_EN_0    <=  '1';
                        Bypass_EN_1    <=  '0';
                        Bypass_EN_2    <=  '0';
                        Bypass_EN_3    <=  '0';
                        Bypass_EN_4    <=  '0';
                        Bypass_EN_5    <=  '0';
                        Bypass_EN_6    <=  '0';
                        Bypass_EN_7    <=  '0';
                        Hold_Ctrl_0    <=  '0';
                        Hold_Ctrl_1    <=  '0';
                        Hold_Ctrl_2    <=  '0';
                        Hold_Ctrl_3    <=  '0';
                        Hold_Ctrl_4    <=  '0';
                        Hold_Ctrl_5    <=  '0';
                        Hold_Ctrl_6    <=  '0';
                        Hold_Ctrl_7    <=  '0';
                        DFF_Ctrl_0     <=  '0';
                        DFF_Ctrl_1     <=  '0';
                        DFF_Ctrl_2     <=  '0';
                        DFF_Ctrl_3     <=  '0';
                        DFF_Ctrl_4     <=  '0';
                        DFF_Ctrl_5     <=  '0';
                        DFF_Ctrl_6     <=  '0';
                        DFF_Ctrl_7     <=  '0';
                        hold_seg_0     <=  '1';
                        hold_seg_1     <=  '1';
                        hold_seg_2     <=  '1';
                        hold_seg_3     <=  '1';
                        hold_seg_4     <=  '1';
                        hold_seg_5     <=  '1';
                        hold_seg_6     <=  '1';
                        hold_seg_7     <=  '0';
                        in_ctrl_all_cb <=  '1';
                        hold_all_out   <=  '0';
                        in_ctrl_all_out<=  '1';
                        counter_en     <=  '0';
                        currentstate   <= state_14;					
                    WHEN state_14		 =>
                        hold_all_in    <=  '0';
                        hold_buf_3     <=  '1';
                        hold_buf_2     <=  '1';
                        hold_buf_1     <=  '1';
                        in_ctrl_buf_3  <=  '0';
                        in_ctrl_buf_2  <=  '0';
                        in_ctrl_buf_1  <=  '0';
                        pos_hold_ctrl  <=  '0';
                        Shuf_Ctrl_1    <=  "000";
                        Shuf_Ctrl_2    <=  "000";
                        Shuf_Ctrl_3    <=  "000";
                        Shuf_Ctrl_4    <=  "000";
                        Shuf_Ctrl_5    <=  "000";
                        Shuf_Ctrl_6    <=  "000";
                        Shuf_Ctrl_7    <=  "000";
                        Shuf_Ctrl_8    <=  "000";
                        Type_Sel_1     <=  "000";
                        Type_Sel_2     <=  "000";
                        Type_Sel_3     <=  "000";
                        Type_Sel_4     <=  "000";
                        Type_Sel_5     <=  "000";
                        Type_Sel_6     <=  "000";
                        Type_Sel_7     <=  "000";
                        Type_Sel_8     <=  "000";
                        Bypass_Sel_0   <=  "000";
                        Bypass_Sel_1   <=  "000";
                        Bypass_Sel_2   <=  "000";
                        Bypass_Sel_3   <=  "000";
                        Bypass_Sel_4   <=  "000";
                        Bypass_Sel_5   <=  "000";
                        Bypass_Sel_6   <=  "000";
                        Bypass_Sel_7   <=  "000";
                        DeShuf_Ctrl_0  <=  "000";
                        DeShuf_Ctrl_1  <=  "000";
                        DeShuf_Ctrl_2  <=  "000";
                        DeShuf_Ctrl_3  <=  "000";
                        DeShuf_Ctrl_4  <=  "000";
                        DeShuf_Ctrl_5  <=  "000";
                        DeShuf_Ctrl_6  <=  "000";
                        DeShuf_Ctrl_7  <=  "000";
                        Bypass_EN_0    <=  '0';
                        Bypass_EN_1    <=  '0';
                        Bypass_EN_2    <=  '0';
                        Bypass_EN_3    <=  '0';
                        Bypass_EN_4    <=  '0';
                        Bypass_EN_5    <=  '0';
                        Bypass_EN_6    <=  '0';
                        Bypass_EN_7    <=  '0';
                        Hold_Ctrl_0    <=  '0';
                        Hold_Ctrl_1    <=  '0';
                        Hold_Ctrl_2    <=  '0';
                        Hold_Ctrl_3    <=  '0';
                        Hold_Ctrl_4    <=  '0';
                        Hold_Ctrl_5    <=  '0';
                        Hold_Ctrl_6    <=  '0';
                        Hold_Ctrl_7    <=  '0';
                        DFF_Ctrl_0     <=  '0';
                        DFF_Ctrl_1     <=  '0';
                        DFF_Ctrl_2     <=  '0';
                        DFF_Ctrl_3     <=  '0';
                        DFF_Ctrl_4     <=  '0';
                        DFF_Ctrl_5     <=  '0';
                        DFF_Ctrl_6     <=  '0';
                        DFF_Ctrl_7     <=  '0';
                        hold_seg_0     <=  '0';
                        hold_seg_1     <=  '0';
                        hold_seg_2     <=  '0';
                        hold_seg_3     <=  '0';
                        hold_seg_4     <=  '0';
                        hold_seg_5     <=  '0';
                        hold_seg_6     <=  '0';
                        hold_seg_7     <=  '0';
                        in_ctrl_all_cb <=  '0';
                        hold_all_out   <=  '0';
                        in_ctrl_all_out<=  '1';
                        counter_en     <=  '1';
                        currentstate   <= state_15;					
                    WHEN state_15		 =>
                        hold_all_in    <=  '0';
                        hold_buf_3     <=  '1';
                        hold_buf_2     <=  '1';
                        hold_buf_1     <=  '1';
                        in_ctrl_buf_3  <=  '0';
                        in_ctrl_buf_2  <=  '0';
                        in_ctrl_buf_1  <=  '0';
                        pos_hold_ctrl  <=  '0';
                        Shuf_Ctrl_1    <=  "000";
                        Shuf_Ctrl_2    <=  "000";
                        Shuf_Ctrl_3    <=  "000";
                        Shuf_Ctrl_4    <=  "000";
                        Shuf_Ctrl_5    <=  "000";
                        Shuf_Ctrl_6    <=  "000";
                        Shuf_Ctrl_7    <=  "000";
                        Shuf_Ctrl_8    <=  "000";
                        Type_Sel_1     <=  "000";
                        Type_Sel_2     <=  "000";
                        Type_Sel_3     <=  "000";
                        Type_Sel_4     <=  "000";
                        Type_Sel_5     <=  "000";
                        Type_Sel_6     <=  "000";
                        Type_Sel_7     <=  "000";
                        Type_Sel_8     <=  "000";
                        Bypass_Sel_0   <=  "000";
                        Bypass_Sel_1   <=  "000";
                        Bypass_Sel_2   <=  "000";
                        Bypass_Sel_3   <=  "000";
                        Bypass_Sel_4   <=  "000";
                        Bypass_Sel_5   <=  "000";
                        Bypass_Sel_6   <=  "000";
                        Bypass_Sel_7   <=  "000";
                        DeShuf_Ctrl_0  <=  "000";
                        DeShuf_Ctrl_1  <=  "000";
                        DeShuf_Ctrl_2  <=  "000";
                        DeShuf_Ctrl_3  <=  "000";
                        DeShuf_Ctrl_4  <=  "000";
                        DeShuf_Ctrl_5  <=  "000";
                        DeShuf_Ctrl_6  <=  "000";
                        DeShuf_Ctrl_7  <=  "000";
                        Bypass_EN_0    <=  '0';
                        Bypass_EN_1    <=  '0';
                        Bypass_EN_2    <=  '0';
                        Bypass_EN_3    <=  '0';
                        Bypass_EN_4    <=  '0';
                        Bypass_EN_5    <=  '0';
                        Bypass_EN_6    <=  '0';
                        Bypass_EN_7    <=  '0';
                        Hold_Ctrl_0    <=  '0';
                        Hold_Ctrl_1    <=  '0';
                        Hold_Ctrl_2    <=  '0';
                        Hold_Ctrl_3    <=  '0';
                        Hold_Ctrl_4    <=  '0';
                        Hold_Ctrl_5    <=  '0';
                        Hold_Ctrl_6    <=  '0';
                        Hold_Ctrl_7    <=  '0';
                        DFF_Ctrl_0     <=  '0';
                        DFF_Ctrl_1     <=  '0';
                        DFF_Ctrl_2     <=  '0';
                        DFF_Ctrl_3     <=  '0';
                        DFF_Ctrl_4     <=  '0';
                        DFF_Ctrl_5     <=  '0';
                        DFF_Ctrl_6     <=  '0';
                        DFF_Ctrl_7     <=  '0';
                        hold_seg_0     <=  '0';
                        hold_seg_1     <=  '0';
                        hold_seg_2     <=  '0';
                        hold_seg_3     <=  '0';
                        hold_seg_4     <=  '0';
                        hold_seg_5     <=  '0';
                        hold_seg_6     <=  '0';
                        hold_seg_7     <=  '0';
                        in_ctrl_all_cb <=  '0';
                        hold_all_out   <=  '0';
                        in_ctrl_all_out<=  '1';
                        counter_en     <=  '0';
                        currentstate   <= state_16;					
                    WHEN state_16		 =>
                        hold_all_in    <=  '0';
                        hold_buf_3     <=  '1';
                        hold_buf_2     <=  '1';
                        hold_buf_1     <=  '1';
                        in_ctrl_buf_3  <=  '0';
                        in_ctrl_buf_2  <=  '0';
                        in_ctrl_buf_1  <=  '0';
                        pos_hold_ctrl  <=  '0';
                        Shuf_Ctrl_1    <=  "000";
                        Shuf_Ctrl_2    <=  "000";
                        Shuf_Ctrl_3    <=  "000";
                        Shuf_Ctrl_4    <=  "000";
                        Shuf_Ctrl_5    <=  "000";
                        Shuf_Ctrl_6    <=  "000";
                        Shuf_Ctrl_7    <=  "000";
                        Shuf_Ctrl_8    <=  "000";
                        Type_Sel_1     <=  "000";
                        Type_Sel_2     <=  "000";
                        Type_Sel_3     <=  "000";
                        Type_Sel_4     <=  "000";
                        Type_Sel_5     <=  "000";
                        Type_Sel_6     <=  "000";
                        Type_Sel_7     <=  "000";
                        Type_Sel_8     <=  "000";
                        Bypass_Sel_0   <=  "000";
                        Bypass_Sel_1   <=  "000";
                        Bypass_Sel_2   <=  "000";
                        Bypass_Sel_3   <=  "000";
                        Bypass_Sel_4   <=  "000";
                        Bypass_Sel_5   <=  "000";
                        Bypass_Sel_6   <=  "000";
                        Bypass_Sel_7   <=  "000";
                        DeShuf_Ctrl_0  <=  "000";
                        DeShuf_Ctrl_1  <=  "000";
                        DeShuf_Ctrl_2  <=  "000";
                        DeShuf_Ctrl_3  <=  "000";
                        DeShuf_Ctrl_4  <=  "000";
                        DeShuf_Ctrl_5  <=  "000";
                        DeShuf_Ctrl_6  <=  "000";
                        DeShuf_Ctrl_7  <=  "000";
                        Bypass_EN_0    <=  '0';
                        Bypass_EN_1    <=  '0';
                        Bypass_EN_2    <=  '0';
                        Bypass_EN_3    <=  '0';
                        Bypass_EN_4    <=  '0';
                        Bypass_EN_5    <=  '0';
                        Bypass_EN_6    <=  '0';
                        Bypass_EN_7    <=  '0';
                        Hold_Ctrl_0    <=  '0';
                        Hold_Ctrl_1    <=  '0';
                        Hold_Ctrl_2    <=  '0';
                        Hold_Ctrl_3    <=  '0';
                        Hold_Ctrl_4    <=  '0';
                        Hold_Ctrl_5    <=  '0';
                        Hold_Ctrl_6    <=  '0';
                        Hold_Ctrl_7    <=  '0';
                        DFF_Ctrl_0     <=  '0';
                        DFF_Ctrl_1     <=  '0';
                        DFF_Ctrl_2     <=  '0';
                        DFF_Ctrl_3     <=  '0';
                        DFF_Ctrl_4     <=  '0';
                        DFF_Ctrl_5     <=  '0';
                        DFF_Ctrl_6     <=  '0';
                        DFF_Ctrl_7     <=  '0';
                        hold_seg_0     <=  '0';
                        hold_seg_1     <=  '0';
                        hold_seg_2     <=  '0';
                        hold_seg_3     <=  '0';
                        hold_seg_4     <=  '0';
                        hold_seg_5     <=  '0';
                        hold_seg_6     <=  '0';
                        hold_seg_7     <=  '0';
                        in_ctrl_all_cb <=  '0';
                        hold_all_out   <=  '0';
                        in_ctrl_all_out<=  '1';
                        counter_en     <=  '0';
                        currentstate   <= state_17;					
                    WHEN state_17		 =>
                        hold_all_in    <=  '0';
                        hold_buf_3     <=  '1';
                        hold_buf_2     <=  '1';
                        hold_buf_1     <=  '1';
                        in_ctrl_buf_3  <=  '0';
                        in_ctrl_buf_2  <=  '0';
                        in_ctrl_buf_1  <=  '0';
                        pos_hold_ctrl  <=  '0';
                        Shuf_Ctrl_1    <=  "000";
                        Shuf_Ctrl_2    <=  "000";
                        Shuf_Ctrl_3    <=  "000";
                        Shuf_Ctrl_4    <=  "000";
                        Shuf_Ctrl_5    <=  "000";
                        Shuf_Ctrl_6    <=  "000";
                        Shuf_Ctrl_7    <=  "000";
                        Shuf_Ctrl_8    <=  "000";
                        Type_Sel_1     <=  "000";
                        Type_Sel_2     <=  "000";
                        Type_Sel_3     <=  "000";
                        Type_Sel_4     <=  "000";
                        Type_Sel_5     <=  "000";
                        Type_Sel_6     <=  "000";
                        Type_Sel_7     <=  "000";
                        Type_Sel_8     <=  "000";
                        Bypass_Sel_0   <=  "000";
                        Bypass_Sel_1   <=  "000";
                        Bypass_Sel_2   <=  "000";
                        Bypass_Sel_3   <=  "000";
                        Bypass_Sel_4   <=  "000";
                        Bypass_Sel_5   <=  "000";
                        Bypass_Sel_6   <=  "000";
                        Bypass_Sel_7   <=  "000";
                        DeShuf_Ctrl_0  <=  "000";
                        DeShuf_Ctrl_1  <=  "000";
                        DeShuf_Ctrl_2  <=  "000";
                        DeShuf_Ctrl_3  <=  "000";
                        DeShuf_Ctrl_4  <=  "000";
                        DeShuf_Ctrl_5  <=  "000";
                        DeShuf_Ctrl_6  <=  "000";
                        DeShuf_Ctrl_7  <=  "000";
                        Bypass_EN_0    <=  '0';
                        Bypass_EN_1    <=  '0';
                        Bypass_EN_2    <=  '0';
                        Bypass_EN_3    <=  '0';
                        Bypass_EN_4    <=  '0';
                        Bypass_EN_5    <=  '0';
                        Bypass_EN_6    <=  '0';
                        Bypass_EN_7    <=  '0';
                        Hold_Ctrl_0    <=  '0';
                        Hold_Ctrl_1    <=  '0';
                        Hold_Ctrl_2    <=  '0';
                        Hold_Ctrl_3    <=  '0';
                        Hold_Ctrl_4    <=  '0';
                        Hold_Ctrl_5    <=  '0';
                        Hold_Ctrl_6    <=  '0';
                        Hold_Ctrl_7    <=  '0';
                        DFF_Ctrl_0     <=  '0';
                        DFF_Ctrl_1     <=  '0';
                        DFF_Ctrl_2     <=  '0';
                        DFF_Ctrl_3     <=  '0';
                        DFF_Ctrl_4     <=  '0';
                        DFF_Ctrl_5     <=  '0';
                        DFF_Ctrl_6     <=  '0';
                        DFF_Ctrl_7     <=  '0';
                        hold_seg_0     <=  '0';
                        hold_seg_1     <=  '0';
                        hold_seg_2     <=  '0';
                        hold_seg_3     <=  '0';
                        hold_seg_4     <=  '0';
                        hold_seg_5     <=  '0';
                        hold_seg_6     <=  '0';
                        hold_seg_7     <=  '0';
                        in_ctrl_all_cb <=  '0';
                        hold_all_out   <=  '0';
                        in_ctrl_all_out<=  '1';
                        counter_en     <=  '0';
                        currentstate   <= state_18;				
                    WHEN state_18		 =>
                        hold_all_in    <=  '0';
                        hold_buf_3     <=  '1';
                        hold_buf_2     <=  '1';
                        hold_buf_1     <=  '1';
                        in_ctrl_buf_3  <=  '0';
                        in_ctrl_buf_2  <=  '0';
                        in_ctrl_buf_1  <=  '0';
                        pos_hold_ctrl  <=  '0';
                        Shuf_Ctrl_1    <=  "000";
                        Shuf_Ctrl_2    <=  "000";
                        Shuf_Ctrl_3    <=  "000";
                        Shuf_Ctrl_4    <=  "000";
                        Shuf_Ctrl_5    <=  "000";
                        Shuf_Ctrl_6    <=  "000";
                        Shuf_Ctrl_7    <=  "000";
                        Shuf_Ctrl_8    <=  "000";
                        Type_Sel_1     <=  "000";
                        Type_Sel_2     <=  "000";
                        Type_Sel_3     <=  "000";
                        Type_Sel_4     <=  "000";
                        Type_Sel_5     <=  "000";
                        Type_Sel_6     <=  "000";
                        Type_Sel_7     <=  "000";
                        Type_Sel_8     <=  "000";
                        Bypass_Sel_0   <=  "000";
                        Bypass_Sel_1   <=  "000";
                        Bypass_Sel_2   <=  "000";
                        Bypass_Sel_3   <=  "000";
                        Bypass_Sel_4   <=  "000";
                        Bypass_Sel_5   <=  "000";
                        Bypass_Sel_6   <=  "000";
                        Bypass_Sel_7   <=  "000";
                        DeShuf_Ctrl_0  <=  "000";
                        DeShuf_Ctrl_1  <=  "000";
                        DeShuf_Ctrl_2  <=  "000";
                        DeShuf_Ctrl_3  <=  "000";
                        DeShuf_Ctrl_4  <=  "000";
                        DeShuf_Ctrl_5  <=  "000";
                        DeShuf_Ctrl_6  <=  "000";
                        DeShuf_Ctrl_7  <=  "000";
                        Bypass_EN_0    <=  '0';
                        Bypass_EN_1    <=  '0';
                        Bypass_EN_2    <=  '0';
                        Bypass_EN_3    <=  '0';
                        Bypass_EN_4    <=  '0';
                        Bypass_EN_5    <=  '0';
                        Bypass_EN_6    <=  '0';
                        Bypass_EN_7    <=  '0';
                        Hold_Ctrl_0    <=  '0';
                        Hold_Ctrl_1    <=  '0';
                        Hold_Ctrl_2    <=  '0';
                        Hold_Ctrl_3    <=  '0';
                        Hold_Ctrl_4    <=  '0';
                        Hold_Ctrl_5    <=  '0';
                        Hold_Ctrl_6    <=  '0';
                        Hold_Ctrl_7    <=  '0';
                        DFF_Ctrl_0     <=  '0';
                        DFF_Ctrl_1     <=  '0';
                        DFF_Ctrl_2     <=  '0';
                        DFF_Ctrl_3     <=  '0';
                        DFF_Ctrl_4     <=  '0';
                        DFF_Ctrl_5     <=  '0';
                        DFF_Ctrl_6     <=  '0';
                        DFF_Ctrl_7     <=  '0';
                        hold_seg_0     <=  '0';
                        hold_seg_1     <=  '0';
                        hold_seg_2     <=  '0';
                        hold_seg_3     <=  '0';
                        hold_seg_4     <=  '0';
                        hold_seg_5     <=  '0';
                        hold_seg_6     <=  '0';
                        hold_seg_7     <=  '0';
                        in_ctrl_all_cb <=  '0';
                        hold_all_out   <=  '0';
                        in_ctrl_all_out<=  '1';
                        counter_en     <=  '0';
                        currentstate   <= state_19;					
                    WHEN state_19		 =>
                        hold_all_in    <=  '0';
                        hold_buf_3     <=  '1';
                        hold_buf_2     <=  '1';
                        hold_buf_1     <=  '1';
                        in_ctrl_buf_3  <=  '0';
                        in_ctrl_buf_2  <=  '0';
                        in_ctrl_buf_1  <=  '0';
                        pos_hold_ctrl  <=  '0';
                        Shuf_Ctrl_1    <=  "000";
                        Shuf_Ctrl_2    <=  "000";
                        Shuf_Ctrl_3    <=  "000";
                        Shuf_Ctrl_4    <=  "000";
                        Shuf_Ctrl_5    <=  "000";
                        Shuf_Ctrl_6    <=  "000";
                        Shuf_Ctrl_7    <=  "000";
                        Shuf_Ctrl_8    <=  "000";
                        Type_Sel_1     <=  "000";
                        Type_Sel_2     <=  "000";
                        Type_Sel_3     <=  "000";
                        Type_Sel_4     <=  "000";
                        Type_Sel_5     <=  "000";
                        Type_Sel_6     <=  "000";
                        Type_Sel_7     <=  "000";
                        Type_Sel_8     <=  "000";
                        Bypass_Sel_0   <=  "000";
                        Bypass_Sel_1   <=  "000";
                        Bypass_Sel_2   <=  "000";
                        Bypass_Sel_3   <=  "000";
                        Bypass_Sel_4   <=  "000";
                        Bypass_Sel_5   <=  "000";
                        Bypass_Sel_6   <=  "000";
                        Bypass_Sel_7   <=  "000";
                        DeShuf_Ctrl_0  <=  "000";
                        DeShuf_Ctrl_1  <=  "000";
                        DeShuf_Ctrl_2  <=  "000";
                        DeShuf_Ctrl_3  <=  "000";
                        DeShuf_Ctrl_4  <=  "000";
                        DeShuf_Ctrl_5  <=  "000";
                        DeShuf_Ctrl_6  <=  "000";
                        DeShuf_Ctrl_7  <=  "000";
                        Bypass_EN_0    <=  '0';
                        Bypass_EN_1    <=  '0';
                        Bypass_EN_2    <=  '0';
                        Bypass_EN_3    <=  '0';
                        Bypass_EN_4    <=  '0';
                        Bypass_EN_5    <=  '0';
                        Bypass_EN_6    <=  '0';
                        Bypass_EN_7    <=  '0';
                        Hold_Ctrl_0    <=  '0';
                        Hold_Ctrl_1    <=  '0';
                        Hold_Ctrl_2    <=  '0';
                        Hold_Ctrl_3    <=  '0';
                        Hold_Ctrl_4    <=  '0';
                        Hold_Ctrl_5    <=  '0';
                        Hold_Ctrl_6    <=  '0';
                        Hold_Ctrl_7    <=  '0';
                        DFF_Ctrl_0     <=  '0';
                        DFF_Ctrl_1     <=  '0';
                        DFF_Ctrl_2     <=  '0';
                        DFF_Ctrl_3     <=  '0';
                        DFF_Ctrl_4     <=  '0';
                        DFF_Ctrl_5     <=  '0';
                        DFF_Ctrl_6     <=  '0';
                        DFF_Ctrl_7     <=  '0';
                        hold_seg_0     <=  '0';
                        hold_seg_1     <=  '0';
                        hold_seg_2     <=  '0';
                        hold_seg_3     <=  '0';
                        hold_seg_4     <=  '0';
                        hold_seg_5     <=  '0';
                        hold_seg_6     <=  '0';
                        hold_seg_7     <=  '0';
                        in_ctrl_all_cb <=  '0';
                        hold_all_out   <=  '0';
                        in_ctrl_all_out<=  '1';
                        counter_en     <=  '0';
                        currentstate   <= state_20;					
                    WHEN state_20		 =>
                        hold_all_in    <=  '0';
                        hold_buf_3     <=  '1';
                        hold_buf_2     <=  '1';
                        hold_buf_1     <=  '1';
                        in_ctrl_buf_3  <=  '0';
                        in_ctrl_buf_2  <=  '0';
                        in_ctrl_buf_1  <=  '0';
                        pos_hold_ctrl  <=  '0';
                        Shuf_Ctrl_1    <=  "000";
                        Shuf_Ctrl_2    <=  "000";
                        Shuf_Ctrl_3    <=  "000";
                        Shuf_Ctrl_4    <=  "000";
                        Shuf_Ctrl_5    <=  "000";
                        Shuf_Ctrl_6    <=  "000";
                        Shuf_Ctrl_7    <=  "000";
                        Shuf_Ctrl_8    <=  "000";
                        Type_Sel_1     <=  "000";
                        Type_Sel_2     <=  "000";
                        Type_Sel_3     <=  "000";
                        Type_Sel_4     <=  "000";
                        Type_Sel_5     <=  "000";
                        Type_Sel_6     <=  "000";
                        Type_Sel_7     <=  "000";
                        Type_Sel_8     <=  "000";
                        Bypass_Sel_0   <=  "000";
                        Bypass_Sel_1   <=  "000";
                        Bypass_Sel_2   <=  "000";
                        Bypass_Sel_3   <=  "000";
                        Bypass_Sel_4   <=  "000";
                        Bypass_Sel_5   <=  "000";
                        Bypass_Sel_6   <=  "000";
                        Bypass_Sel_7   <=  "000";
                        DeShuf_Ctrl_0  <=  "000";
                        DeShuf_Ctrl_1  <=  "000";
                        DeShuf_Ctrl_2  <=  "000";
                        DeShuf_Ctrl_3  <=  "000";
                        DeShuf_Ctrl_4  <=  "000";
                        DeShuf_Ctrl_5  <=  "000";
                        DeShuf_Ctrl_6  <=  "000";
                        DeShuf_Ctrl_7  <=  "000";
                        Bypass_EN_0    <=  '0';
                        Bypass_EN_1    <=  '0';
                        Bypass_EN_2    <=  '0';
                        Bypass_EN_3    <=  '0';
                        Bypass_EN_4    <=  '0';
                        Bypass_EN_5    <=  '0';
                        Bypass_EN_6    <=  '0';
                        Bypass_EN_7    <=  '0';
                        Hold_Ctrl_0    <=  '0';
                        Hold_Ctrl_1    <=  '0';
                        Hold_Ctrl_2    <=  '0';
                        Hold_Ctrl_3    <=  '0';
                        Hold_Ctrl_4    <=  '0';
                        Hold_Ctrl_5    <=  '0';
                        Hold_Ctrl_6    <=  '0';
                        Hold_Ctrl_7    <=  '0';
                        DFF_Ctrl_0     <=  '0';
                        DFF_Ctrl_1     <=  '0';
                        DFF_Ctrl_2     <=  '0';
                        DFF_Ctrl_3     <=  '0';
                        DFF_Ctrl_4     <=  '0';
                        DFF_Ctrl_5     <=  '0';
                        DFF_Ctrl_6     <=  '0';
                        DFF_Ctrl_7     <=  '0';
                        hold_seg_0     <=  '0';
                        hold_seg_1     <=  '0';
                        hold_seg_2     <=  '0';
                        hold_seg_3     <=  '0';
                        hold_seg_4     <=  '0';
                        hold_seg_5     <=  '0';
                        hold_seg_6     <=  '0';
                        hold_seg_7     <=  '0';
                        in_ctrl_all_cb <=  '0';
                        hold_all_out   <=  '0';
                        in_ctrl_all_out<=  '1';
                        counter_en     <=  '0';
                        currentstate   <= state_21;					
                    WHEN state_21		 =>		
                        hold_all_in    <=  '0';
                        hold_buf_3     <=  '1';
                        hold_buf_2     <=  '1';
                        hold_buf_1     <=  '1';
                        in_ctrl_buf_3  <=  '0';
                        in_ctrl_buf_2  <=  '0';
                        in_ctrl_buf_1  <=  '0';
                        pos_hold_ctrl  <=  '0';
                        Shuf_Ctrl_1    <=  "000";
                        Shuf_Ctrl_2    <=  "000";
                        Shuf_Ctrl_3    <=  "000";
                        Shuf_Ctrl_4    <=  "000";
                        Shuf_Ctrl_5    <=  "000";
                        Shuf_Ctrl_6    <=  "000";
                        Shuf_Ctrl_7    <=  "000";
                        Shuf_Ctrl_8    <=  "000";
                        Type_Sel_1     <=  "000";
                        Type_Sel_2     <=  "000";
                        Type_Sel_3     <=  "000";
                        Type_Sel_4     <=  "000";
                        Type_Sel_5     <=  "000";
                        Type_Sel_6     <=  "000";
                        Type_Sel_7     <=  "000";
                        Type_Sel_8     <=  "000";
                        Bypass_Sel_0   <=  "000";
                        Bypass_Sel_1   <=  "000";
                        Bypass_Sel_2   <=  "000";
                        Bypass_Sel_3   <=  "000";
                        Bypass_Sel_4   <=  "000";
                        Bypass_Sel_5   <=  "000";
                        Bypass_Sel_6   <=  "000";
                        Bypass_Sel_7   <=  "000";
                        DeShuf_Ctrl_0  <=  "000";
                        DeShuf_Ctrl_1  <=  "000";
                        DeShuf_Ctrl_2  <=  "000";
                        DeShuf_Ctrl_3  <=  "000";
                        DeShuf_Ctrl_4  <=  "000";
                        DeShuf_Ctrl_5  <=  "000";
                        DeShuf_Ctrl_6  <=  "000";
                        DeShuf_Ctrl_7  <=  "000";
                        Bypass_EN_0    <=  '0';
                        Bypass_EN_1    <=  '0';
                        Bypass_EN_2    <=  '0';
                        Bypass_EN_3    <=  '0';
                        Bypass_EN_4    <=  '0';
                        Bypass_EN_5    <=  '0';
                        Bypass_EN_6    <=  '0';
                        Bypass_EN_7    <=  '0';
                        Hold_Ctrl_0    <=  '0';
                        Hold_Ctrl_1    <=  '0';
                        Hold_Ctrl_2    <=  '0';
                        Hold_Ctrl_3    <=  '0';
                        Hold_Ctrl_4    <=  '0';
                        Hold_Ctrl_5    <=  '0';
                        Hold_Ctrl_6    <=  '0';
                        Hold_Ctrl_7    <=  '0';
                        DFF_Ctrl_0     <=  '0';
                        DFF_Ctrl_1     <=  '0';
                        DFF_Ctrl_2     <=  '0';
                        DFF_Ctrl_3     <=  '0';
                        DFF_Ctrl_4     <=  '0';
                        DFF_Ctrl_5     <=  '0';
                        DFF_Ctrl_6     <=  '0';
                        DFF_Ctrl_7     <=  '0';
                        hold_seg_0     <=  '0';
                        hold_seg_1     <=  '0';
                        hold_seg_2     <=  '0';
                        hold_seg_3     <=  '0';
                        hold_seg_4     <=  '0';
                        hold_seg_5     <=  '0';
                        hold_seg_6     <=  '0';
                        hold_seg_7     <=  '0';
                        in_ctrl_all_cb <=  '0';
                        hold_all_out   <=  '0';
                        in_ctrl_all_out<=  '0';
                        counter_en     <=  '0';
                        currentstate   <= state_22;
					WHEN state_22		 =>		
                        hold_all_in    <=  '0';
                        hold_buf_3     <=  '1';
                        hold_buf_2     <=  '1';
                        hold_buf_1     <=  '1';
                        in_ctrl_buf_3  <=  '0';
                        in_ctrl_buf_2  <=  '0';
                        in_ctrl_buf_1  <=  '0';
                        pos_hold_ctrl  <=  '0';
                        Shuf_Ctrl_1    <=  "000";
                        Shuf_Ctrl_2    <=  "000";
                        Shuf_Ctrl_3    <=  "000";
                        Shuf_Ctrl_4    <=  "000";
                        Shuf_Ctrl_5    <=  "000";
                        Shuf_Ctrl_6    <=  "000";
                        Shuf_Ctrl_7    <=  "000";
                        Shuf_Ctrl_8    <=  "000";
                        Type_Sel_1     <=  "000";
                        Type_Sel_2     <=  "000";
                        Type_Sel_3     <=  "000";
                        Type_Sel_4     <=  "000";
                        Type_Sel_5     <=  "000";
                        Type_Sel_6     <=  "000";
                        Type_Sel_7     <=  "000";
                        Type_Sel_8     <=  "000";
                        Bypass_Sel_0   <=  "000";
                        Bypass_Sel_1   <=  "000";
                        Bypass_Sel_2   <=  "000";
                        Bypass_Sel_3   <=  "000";
                        Bypass_Sel_4   <=  "000";
                        Bypass_Sel_5   <=  "000";
                        Bypass_Sel_6   <=  "000";
                        Bypass_Sel_7   <=  "000";
                        DeShuf_Ctrl_0  <=  "000";
                        DeShuf_Ctrl_1  <=  "000";
                        DeShuf_Ctrl_2  <=  "000";
                        DeShuf_Ctrl_3  <=  "000";
                        DeShuf_Ctrl_4  <=  "000";
                        DeShuf_Ctrl_5  <=  "000";
                        DeShuf_Ctrl_6  <=  "000";
                        DeShuf_Ctrl_7  <=  "000";
                        Bypass_EN_0    <=  '0';
                        Bypass_EN_1    <=  '0';
                        Bypass_EN_2    <=  '0';
                        Bypass_EN_3    <=  '0';
                        Bypass_EN_4    <=  '0';
                        Bypass_EN_5    <=  '0';
                        Bypass_EN_6    <=  '0';
                        Bypass_EN_7    <=  '0';
                        Hold_Ctrl_0    <=  '0';
                        Hold_Ctrl_1    <=  '0';
                        Hold_Ctrl_2    <=  '0';
                        Hold_Ctrl_3    <=  '0';
                        Hold_Ctrl_4    <=  '0';
                        Hold_Ctrl_5    <=  '0';
                        Hold_Ctrl_6    <=  '0';
                        Hold_Ctrl_7    <=  '0';
                        DFF_Ctrl_0     <=  '0';
                        DFF_Ctrl_1     <=  '0';
                        DFF_Ctrl_2     <=  '0';
                        DFF_Ctrl_3     <=  '0';
                        DFF_Ctrl_4     <=  '0';
                        DFF_Ctrl_5     <=  '0';
                        DFF_Ctrl_6     <=  '0';
                        DFF_Ctrl_7     <=  '0';
                        hold_seg_0     <=  '1';
                        hold_seg_1     <=  '1';
                        hold_seg_2     <=  '1';
                        hold_seg_3     <=  '1';
                        hold_seg_4     <=  '1';
                        hold_seg_5     <=  '1';
                        hold_seg_6     <=  '1';
                        hold_seg_7     <=  '1';
                        in_ctrl_all_cb <=  '1';
                        hold_all_out   <=  '0';
                        in_ctrl_all_out<=  '0';
                        counter_en     <=  '0';
                        currentstate   <= state_0;					
				END CASE;
			ELSE
				currentstate <= currentstate;
			END IF;
		END IF;		
	END PROCESS;
END behavioral;
